// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 15:54:18 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3,
    i4  );
  input  i0, i1, i2, i3;
  output i4;
  assign i4 = 1'b1;
endmodule


