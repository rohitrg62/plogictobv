// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:26:57 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8, i9, i10, i11  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8, i9, i10, i11;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
    n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
    n41, n42, n43, n44, n45, n47, n48, n49, n50, n51, n52, n53, n54, n55,
    n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260;
  assign n13 = i0 & i1;
  assign n14 = i3 & n13;
  assign n15 = ~i4 & n14;
  assign n16 = i5 & n15;
  assign n17 = i6 & n16;
  assign n18 = i7 & n17;
  assign n19 = ~i0 & i1;
  assign n20 = i3 & n19;
  assign n21 = i4 & n20;
  assign n22 = ~i5 & n21;
  assign n23 = i6 & n22;
  assign n24 = i7 & n23;
  assign n25 = i6 & n15;
  assign n26 = i7 & n25;
  assign n27 = i4 & n14;
  assign n28 = ~i5 & n27;
  assign n29 = i6 & n28;
  assign n30 = i7 & n29;
  assign n31 = ~i1 & ~i2;
  assign n32 = ~i1 & i2;
  assign n33 = ~i0 & n32;
  assign n34 = ~n31 & ~n33;
  assign n35 = i0 & n32;
  assign n36 = ~i6 & n35;
  assign n37 = n34 & ~n36;
  assign n38 = i6 & n35;
  assign n39 = i4 & n38;
  assign n40 = i7 & n39;
  assign n41 = n37 & ~n40;
  assign n42 = ~i1 & n41;
  assign n43 = ~n18 & ~n42;
  assign n44 = ~n24 & n43;
  assign n45 = ~n26 & n44;
  assign i10 = ~n30 & n45;
  assign n47 = i0 & ~i1;
  assign n48 = i2 & n47;
  assign n49 = i3 & n48;
  assign n50 = ~i6 & n49;
  assign n51 = i7 & n50;
  assign n52 = i10 & n51;
  assign n53 = ~i0 & ~i1;
  assign n54 = i2 & n53;
  assign n55 = i3 & n54;
  assign n56 = i6 & n55;
  assign n57 = ~i7 & n56;
  assign n58 = ~i2 & n47;
  assign n59 = i3 & n58;
  assign n60 = i4 & n59;
  assign n61 = i6 & n60;
  assign n62 = ~i7 & n61;
  assign n63 = i10 & n62;
  assign n64 = ~i0 & ~i2;
  assign n65 = ~i0 & i2;
  assign n66 = ~i3 & n65;
  assign n67 = ~n64 & ~n66;
  assign n68 = i3 & n65;
  assign n69 = n67 & ~n68;
  assign n70 = i0 & ~i6;
  assign n71 = n69 & ~n70;
  assign n72 = i0 & i6;
  assign n73 = ~i1 & n72;
  assign n74 = ~i3 & n73;
  assign n75 = n71 & ~n74;
  assign n76 = i3 & n73;
  assign n77 = ~i7 & n76;
  assign n78 = n75 & ~n77;
  assign n79 = ~n52 & ~n78;
  assign n80 = ~n57 & n79;
  assign i11 = ~n63 & n80;
  assign n82 = ~i2 & n13;
  assign n83 = ~i3 & n82;
  assign n84 = i6 & n83;
  assign n85 = ~i7 & n84;
  assign n86 = i10 & n85;
  assign n87 = ~i11 & n86;
  assign n88 = ~i2 & n19;
  assign n89 = i3 & n88;
  assign n90 = ~i5 & n89;
  assign n91 = i6 & n90;
  assign n92 = ~i10 & n91;
  assign n93 = i11 & n92;
  assign n94 = ~i4 & n89;
  assign n95 = i6 & n94;
  assign n96 = i7 & n95;
  assign n97 = i10 & n96;
  assign n98 = i11 & n97;
  assign n99 = ~i4 & n83;
  assign n100 = i6 & n99;
  assign n101 = i10 & n100;
  assign n102 = ~i11 & n101;
  assign n103 = i3 & n82;
  assign n104 = i4 & n103;
  assign n105 = i5 & n104;
  assign n106 = i6 & n105;
  assign n107 = ~i7 & n106;
  assign n108 = i10 & n107;
  assign n109 = ~i11 & n108;
  assign n110 = i2 & n13;
  assign n111 = i3 & n110;
  assign n112 = ~i4 & n111;
  assign n113 = i6 & n112;
  assign n114 = i7 & n113;
  assign n115 = ~i10 & n114;
  assign n116 = ~i11 & n115;
  assign n117 = i4 & n89;
  assign n118 = i5 & n117;
  assign n119 = i6 & n118;
  assign n120 = ~i7 & n119;
  assign n121 = i10 & n120;
  assign n122 = i11 & n121;
  assign n123 = i5 & n111;
  assign n124 = ~i6 & n123;
  assign n125 = i7 & n124;
  assign n126 = i10 & n125;
  assign n127 = i11 & n126;
  assign n128 = ~i5 & n83;
  assign n129 = i6 & n128;
  assign n130 = i10 & n129;
  assign n131 = ~i11 & n130;
  assign n132 = i2 & n19;
  assign n133 = ~i3 & n132;
  assign n134 = i4 & n133;
  assign n135 = ~i5 & n134;
  assign n136 = i6 & n135;
  assign n137 = i7 & n136;
  assign n138 = i1 & i2;
  assign n139 = i3 & n138;
  assign n140 = ~i5 & n139;
  assign n141 = i6 & n140;
  assign n142 = i7 & n141;
  assign n143 = ~i10 & n142;
  assign n144 = ~i11 & n143;
  assign n145 = ~i4 & n20;
  assign n146 = i6 & n145;
  assign n147 = i7 & n146;
  assign n148 = i10 & n147;
  assign n149 = i11 & n148;
  assign n150 = ~i6 & n111;
  assign n151 = i7 & n150;
  assign n152 = i10 & n151;
  assign n153 = i11 & n152;
  assign n154 = i3 & n132;
  assign n155 = i4 & n154;
  assign n156 = ~i6 & n155;
  assign n157 = i7 & n156;
  assign n158 = i10 & n157;
  assign n159 = i11 & n158;
  assign n160 = i1 & ~i2;
  assign n161 = i1 & ~n160;
  assign n162 = ~i7 & n138;
  assign n163 = ~i6 & n162;
  assign n164 = ~i11 & n163;
  assign n165 = n161 & ~n164;
  assign n166 = i6 & n162;
  assign n167 = ~i10 & n166;
  assign n168 = ~i4 & n167;
  assign n169 = n165 & ~n168;
  assign n170 = i7 & n138;
  assign n171 = n169 & ~n170;
  assign n172 = ~n87 & ~n171;
  assign n173 = ~n93 & n172;
  assign n174 = ~n98 & n173;
  assign n175 = ~n102 & n174;
  assign n176 = ~n109 & n175;
  assign n177 = ~n116 & n176;
  assign n178 = ~n122 & n177;
  assign n179 = ~n127 & n178;
  assign n180 = ~n131 & n179;
  assign n181 = ~n137 & n180;
  assign n182 = ~n144 & n181;
  assign n183 = ~n149 & n182;
  assign n184 = ~n153 & n183;
  assign i8 = ~n159 & n184;
  assign n186 = i0 & i2;
  assign n187 = ~i3 & n186;
  assign n188 = i6 & n187;
  assign n189 = ~i7 & n188;
  assign n190 = ~i8 & n189;
  assign n191 = i10 & n190;
  assign n192 = ~i11 & n191;
  assign n193 = ~i4 & n133;
  assign n194 = i6 & n193;
  assign n195 = i8 & n194;
  assign n196 = i5 & n134;
  assign n197 = ~i6 & n196;
  assign n198 = i7 & n197;
  assign n199 = i8 & n198;
  assign n200 = i1 & i3;
  assign n201 = i4 & n200;
  assign n202 = i5 & n201;
  assign n203 = i6 & n202;
  assign n204 = ~i7 & n203;
  assign n205 = i10 & n204;
  assign n206 = ~i11 & n205;
  assign n207 = ~i3 & n48;
  assign n208 = i4 & n207;
  assign n209 = ~i6 & n208;
  assign n210 = i7 & n209;
  assign n211 = i10 & n210;
  assign n212 = ~i3 & n110;
  assign n213 = i5 & n212;
  assign n214 = ~i6 & n213;
  assign n215 = i7 & n214;
  assign n216 = i8 & n215;
  assign n217 = i10 & n216;
  assign n218 = i11 & n217;
  assign n219 = i4 & n49;
  assign n220 = ~i6 & n219;
  assign n221 = i10 & n220;
  assign n222 = i11 & n221;
  assign n223 = i3 & n47;
  assign n224 = i4 & n223;
  assign n225 = i6 & n224;
  assign n226 = ~i7 & n225;
  assign n227 = i11 & n226;
  assign n228 = ~i6 & n55;
  assign n229 = i7 & n228;
  assign n230 = i11 & n229;
  assign n231 = i7 & n220;
  assign n232 = i10 & n231;
  assign n233 = ~i11 & n232;
  assign n234 = i5 & n21;
  assign n235 = i6 & n234;
  assign n236 = ~i7 & n235;
  assign n237 = i10 & n236;
  assign n238 = i4 & n212;
  assign n239 = ~i6 & n238;
  assign n240 = i7 & n239;
  assign n241 = i8 & n240;
  assign n242 = i10 & n241;
  assign n243 = i11 & n242;
  assign n244 = ~i6 & n154;
  assign n245 = i7 & n244;
  assign n246 = i8 & n245;
  assign n247 = i10 & n246;
  assign n248 = i11 & n247;
  assign n249 = ~n192 & ~n195;
  assign n250 = ~n199 & n249;
  assign n251 = ~n148 & n250;
  assign n252 = ~n206 & n251;
  assign n253 = ~n211 & n252;
  assign n254 = ~n218 & n253;
  assign n255 = ~n222 & n254;
  assign n256 = ~n227 & n255;
  assign n257 = ~n230 & n256;
  assign n258 = ~n233 & n257;
  assign n259 = ~n237 & n258;
  assign n260 = ~n243 & n259;
  assign i9 = ~n248 & n260;
endmodule


