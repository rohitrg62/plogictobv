// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:26:45 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8, i9, i10, i11  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8, i9, i10, i11;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
    n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
    n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
    n55, n56, n57, n58, n59, n60, n61, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
    n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
    n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
    n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
    n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
    n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n369, n370;
  assign n13 = i0 & ~i1;
  assign n14 = ~i2 & n13;
  assign n15 = ~i3 & n14;
  assign n16 = i4 & n15;
  assign n17 = i5 & n16;
  assign n18 = ~i6 & n17;
  assign n19 = i7 & n18;
  assign n20 = ~i4 & n15;
  assign n21 = i5 & n20;
  assign n22 = i6 & n21;
  assign n23 = i7 & n22;
  assign n24 = i0 & ~i2;
  assign n25 = ~i4 & n24;
  assign n26 = i5 & n25;
  assign n27 = ~i6 & n26;
  assign n28 = ~i7 & n27;
  assign n29 = ~i3 & n24;
  assign n30 = i4 & n29;
  assign n31 = i5 & n30;
  assign n32 = i6 & n31;
  assign n33 = ~i7 & n32;
  assign n34 = ~i0 & i1;
  assign n35 = ~i2 & n34;
  assign n36 = ~i3 & n35;
  assign n37 = ~i4 & n36;
  assign n38 = i5 & n37;
  assign n39 = i5 & n36;
  assign n40 = ~i7 & n39;
  assign n41 = ~i0 & ~i1;
  assign n42 = i2 & n41;
  assign n43 = ~i3 & n42;
  assign n44 = ~i4 & n43;
  assign n45 = i5 & n44;
  assign n46 = ~i6 & n45;
  assign n47 = ~i7 & n46;
  assign n48 = ~i6 & n39;
  assign n49 = ~i2 & i3;
  assign n50 = ~i4 & n49;
  assign n51 = i5 & n50;
  assign n52 = ~i6 & n51;
  assign n53 = ~i7 & n52;
  assign n54 = ~n19 & ~n23;
  assign n55 = ~n28 & n54;
  assign n56 = ~n33 & n55;
  assign n57 = ~n38 & n56;
  assign n58 = ~n40 & n57;
  assign n59 = ~n47 & n58;
  assign n60 = ~n48 & n59;
  assign n61 = ~n39 & n60;
  assign i9 = ~n53 & n61;
  assign n63 = i1 & ~i2;
  assign n64 = ~i3 & n63;
  assign n65 = ~i4 & n64;
  assign n66 = ~i5 & n65;
  assign n67 = i7 & n66;
  assign n68 = ~i4 & n63;
  assign n69 = ~i5 & n68;
  assign n70 = i6 & n69;
  assign n71 = ~i7 & n70;
  assign n72 = ~i6 & n31;
  assign n73 = i7 & n72;
  assign n74 = i9 & n73;
  assign n75 = ~i5 & n50;
  assign n76 = i6 & n75;
  assign n77 = ~i7 & n76;
  assign n78 = ~i5 & n25;
  assign n79 = i6 & n78;
  assign n80 = ~i7 & n79;
  assign n81 = ~i2 & n41;
  assign n82 = i3 & n81;
  assign n83 = ~i4 & n82;
  assign n84 = ~i5 & n83;
  assign n85 = i7 & n84;
  assign n86 = ~i4 & n29;
  assign n87 = ~i5 & n86;
  assign n88 = i7 & n87;
  assign n89 = ~i5 & n16;
  assign n90 = i4 & n14;
  assign n91 = i5 & n90;
  assign n92 = ~i6 & n91;
  assign n93 = i7 & n92;
  assign n94 = i9 & n93;
  assign n95 = i4 & n36;
  assign n96 = ~i0 & i2;
  assign n97 = ~i3 & n96;
  assign n98 = ~i4 & n97;
  assign n99 = i5 & n98;
  assign n100 = ~i6 & n99;
  assign n101 = ~i7 & n100;
  assign n102 = i9 & n101;
  assign n103 = ~i5 & n44;
  assign n104 = i6 & n103;
  assign n105 = ~i7 & n104;
  assign n106 = i4 & n35;
  assign n107 = i5 & n106;
  assign n108 = ~i6 & n107;
  assign n109 = i7 & n108;
  assign n110 = i9 & n109;
  assign n111 = i4 & n82;
  assign n112 = i5 & n111;
  assign n113 = ~i6 & n112;
  assign n114 = i7 & n113;
  assign n115 = i9 & n114;
  assign n116 = i5 & n86;
  assign n117 = i6 & n116;
  assign n118 = i7 & n117;
  assign n119 = i9 & n118;
  assign n120 = i4 & n43;
  assign n121 = i5 & n120;
  assign n122 = ~i6 & n121;
  assign n123 = i7 & n122;
  assign n124 = i9 & n123;
  assign n125 = i4 & n97;
  assign n126 = i5 & n125;
  assign n127 = ~i6 & n126;
  assign n128 = i7 & n127;
  assign n129 = i9 & n128;
  assign n130 = i4 & n24;
  assign n131 = i5 & n130;
  assign n132 = ~i6 & n131;
  assign n133 = i7 & n132;
  assign n134 = i9 & n133;
  assign n135 = ~i1 & ~i9;
  assign n136 = ~i1 & i9;
  assign n137 = ~n135 & ~n136;
  assign n138 = ~i1 & n137;
  assign n139 = ~n67 & ~n138;
  assign n140 = ~n71 & n139;
  assign n141 = ~n74 & n140;
  assign n142 = ~n39 & n141;
  assign n143 = ~n77 & n142;
  assign n144 = ~n80 & n143;
  assign n145 = ~n85 & n144;
  assign n146 = ~n88 & n145;
  assign n147 = ~n89 & n146;
  assign n148 = ~n94 & n147;
  assign n149 = ~n95 & n148;
  assign n150 = ~n102 & n149;
  assign n151 = ~n105 & n150;
  assign n152 = ~n110 & n151;
  assign n153 = ~n115 & n152;
  assign n154 = ~n119 & n153;
  assign n155 = ~n124 & n154;
  assign n156 = ~n129 & n155;
  assign i10 = ~n134 & n156;
  assign n158 = i7 & n69;
  assign n159 = ~i10 & n158;
  assign n160 = i5 & n68;
  assign n161 = ~i6 & n160;
  assign n162 = i7 & n161;
  assign n163 = i9 & n162;
  assign n164 = i10 & n163;
  assign n165 = ~i4 & n14;
  assign n166 = i5 & n165;
  assign n167 = ~i6 & n166;
  assign n168 = i7 & n167;
  assign n169 = i9 & n168;
  assign n170 = i10 & n169;
  assign n171 = ~i6 & n78;
  assign n172 = i7 & n171;
  assign n173 = ~i6 & n69;
  assign n174 = i7 & n173;
  assign n175 = i7 & n75;
  assign n176 = ~i10 & n175;
  assign n177 = i7 & n78;
  assign n178 = ~i10 & n177;
  assign n179 = ~i5 & n30;
  assign n180 = ~i10 & n179;
  assign n181 = i4 & n64;
  assign n182 = ~i5 & n181;
  assign n183 = ~i10 & n182;
  assign n184 = n116 & i10;
  assign n185 = i2 & ~i3;
  assign n186 = ~i4 & n185;
  assign n187 = i5 & n186;
  assign n188 = ~i6 & n187;
  assign n189 = ~i7 & n188;
  assign n190 = i9 & n189;
  assign n191 = i10 & n190;
  assign n192 = ~i5 & n111;
  assign n193 = ~i7 & n192;
  assign n194 = i6 & n112;
  assign n195 = ~i7 & n194;
  assign n196 = i9 & n195;
  assign n197 = i10 & n196;
  assign n198 = i5 & n83;
  assign n199 = ~i6 & n198;
  assign n200 = i7 & n199;
  assign n201 = i9 & n200;
  assign n202 = i10 & n201;
  assign n203 = i6 & n107;
  assign n204 = ~i7 & n203;
  assign n205 = i9 & n204;
  assign n206 = i10 & n205;
  assign n207 = ~i7 & n179;
  assign n208 = ~i5 & n186;
  assign n209 = ~i6 & n208;
  assign n210 = i7 & n209;
  assign n211 = i10 & n210;
  assign n212 = ~i5 & n90;
  assign n213 = ~i7 & n212;
  assign n214 = i10 & n213;
  assign n215 = ~i4 & n42;
  assign n216 = ~i5 & n215;
  assign n217 = ~i6 & n216;
  assign n218 = i7 & n217;
  assign n219 = i10 & n218;
  assign n220 = n26 & i9;
  assign n221 = ~i10 & n220;
  assign n222 = ~i5 & n106;
  assign n223 = ~i7 & n222;
  assign n224 = i10 & n223;
  assign n225 = ~n159 & ~n164;
  assign n226 = ~n21 & n225;
  assign n227 = ~n170 & n226;
  assign n228 = ~n39 & n227;
  assign n229 = ~n172 & n228;
  assign n230 = ~n174 & n229;
  assign n231 = ~n176 & n230;
  assign n232 = ~n178 & n231;
  assign n233 = ~n180 & n232;
  assign n234 = ~n183 & n233;
  assign n235 = ~n184 & n234;
  assign n236 = ~n102 & n235;
  assign n237 = ~n191 & n236;
  assign n238 = ~n193 & n237;
  assign n239 = ~n197 & n238;
  assign n240 = ~n202 & n239;
  assign n241 = ~n206 & n240;
  assign n242 = ~n207 & n241;
  assign n243 = ~n211 & n242;
  assign n244 = ~n214 & n243;
  assign n245 = ~n219 & n244;
  assign n246 = ~n221 & ~n245;
  assign i11 = ~n224 & ~n246;
  assign n248 = i5 & n65;
  assign n249 = ~i10 & n248;
  assign n250 = i5 & n64;
  assign n251 = ~i7 & n250;
  assign n252 = ~i11 & n251;
  assign n253 = ~i1 & i2;
  assign n254 = ~i3 & n253;
  assign n255 = i4 & n254;
  assign n256 = ~i5 & n255;
  assign n257 = i6 & n256;
  assign n258 = i7 & n257;
  assign n259 = i10 & n258;
  assign n260 = i11 & n259;
  assign n261 = i4 & n185;
  assign n262 = ~i5 & n261;
  assign n263 = ~i6 & n262;
  assign n264 = ~i7 & n263;
  assign n265 = i11 & n264;
  assign n266 = i4 & n63;
  assign n267 = ~i5 & n266;
  assign n268 = ~i6 & n267;
  assign n269 = ~i7 & n268;
  assign n270 = ~i11 & n269;
  assign n271 = ~i10 & n250;
  assign n272 = ~i11 & n271;
  assign n273 = i4 & n42;
  assign n274 = ~i5 & n273;
  assign n275 = i6 & n274;
  assign n276 = ~i7 & n275;
  assign n277 = i10 & n276;
  assign n278 = i11 & n277;
  assign n279 = i7 & n46;
  assign n280 = i9 & n279;
  assign n281 = i10 & n280;
  assign n282 = i11 & n281;
  assign n283 = ~i10 & n268;
  assign n284 = ~i11 & n283;
  assign n285 = ~i5 & n130;
  assign n286 = ~i6 & n285;
  assign n287 = ~i7 & n286;
  assign n288 = ~i11 & n287;
  assign n289 = ~i10 & n286;
  assign n290 = ~i11 & n289;
  assign n291 = i4 & n96;
  assign n292 = ~i5 & n291;
  assign n293 = ~i6 & n292;
  assign n294 = ~i7 & n293;
  assign n295 = i10 & n294;
  assign n296 = i11 & n295;
  assign n297 = i7 & n188;
  assign n298 = i9 & n297;
  assign n299 = i10 & n298;
  assign n300 = i11 & n299;
  assign n301 = n116 & ~i10;
  assign n302 = i6 & n121;
  assign n303 = ~i7 & n302;
  assign n304 = i9 & n303;
  assign n305 = i10 & n304;
  assign n306 = i11 & n305;
  assign n307 = i6 & n131;
  assign n308 = ~i7 & n307;
  assign n309 = i9 & n308;
  assign n310 = i10 & n309;
  assign n311 = i11 & n310;
  assign n312 = i6 & n126;
  assign n313 = ~i7 & n312;
  assign n314 = i9 & n313;
  assign n315 = i10 & n314;
  assign n316 = i11 & n315;
  assign n317 = ~i5 & n125;
  assign n318 = ~i6 & n317;
  assign n319 = i7 & n318;
  assign n320 = i10 & n319;
  assign n321 = i11 & n320;
  assign n322 = i4 & n253;
  assign n323 = ~i5 & n322;
  assign n324 = i6 & n323;
  assign n325 = ~i7 & n324;
  assign n326 = i10 & n325;
  assign n327 = i11 & n326;
  assign n328 = ~i4 & ~i5;
  assign n329 = i4 & ~i5;
  assign n330 = ~i2 & n329;
  assign n331 = ~i6 & n330;
  assign n332 = ~i10 & n331;
  assign n333 = ~n328 & ~n332;
  assign n334 = i6 & n330;
  assign n335 = i10 & n334;
  assign n336 = ~i3 & n335;
  assign n337 = i0 & n336;
  assign n338 = n333 & ~n337;
  assign n339 = i3 & n335;
  assign n340 = n338 & ~n339;
  assign n341 = i2 & n329;
  assign n342 = ~i1 & n341;
  assign n343 = ~i11 & n342;
  assign n344 = n340 & ~n343;
  assign n345 = i1 & n341;
  assign n346 = n344 & ~n345;
  assign n347 = i5 & ~i7;
  assign n348 = ~i10 & n347;
  assign n349 = n346 & ~n348;
  assign n350 = i5 & i7;
  assign n351 = n349 & ~n350;
  assign n352 = ~n249 & ~n351;
  assign n353 = ~n252 & n352;
  assign n354 = ~n260 & ~n353;
  assign n355 = ~n265 & ~n354;
  assign n356 = ~n270 & n355;
  assign n357 = ~n272 & n356;
  assign n358 = ~n278 & ~n357;
  assign n359 = ~n190 & ~n358;
  assign n360 = ~n282 & n359;
  assign n361 = ~n284 & n360;
  assign n362 = ~n288 & n361;
  assign n363 = ~n290 & n362;
  assign n364 = ~n296 & n363;
  assign n365 = ~n300 & n364;
  assign n366 = ~n301 & n365;
  assign n367 = ~n306 & ~n366;
  assign n368 = ~n311 & n367;
  assign n369 = ~n316 & n368;
  assign n370 = ~n321 & ~n369;
  assign i8 = n327 | n370;
endmodule


