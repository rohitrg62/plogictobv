// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:27:16 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8, i9, i10, i11  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8, i9, i10, i11;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
    n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
    n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
    n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
    n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
    n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
    n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
    n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
    n121, n122, n123, n125, n126, n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
    n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
    n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
    n182, n183, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
    n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
    n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
    n376;
  assign n13 = ~i0 & ~i2;
  assign n14 = ~i4 & n13;
  assign n15 = ~i5 & n14;
  assign n16 = ~i6 & n15;
  assign n17 = ~i7 & n16;
  assign n18 = ~i1 & ~i2;
  assign n19 = ~i4 & n18;
  assign n20 = ~i5 & n19;
  assign n21 = ~i6 & n20;
  assign n22 = ~i7 & n21;
  assign n23 = ~i2 & ~i3;
  assign n24 = ~i4 & n23;
  assign n25 = ~i5 & n24;
  assign n26 = ~i6 & n25;
  assign n27 = ~i7 & n26;
  assign n28 = i3 & n13;
  assign n29 = ~i4 & n28;
  assign n30 = ~i5 & n29;
  assign n31 = ~i6 & n30;
  assign n32 = i7 & n31;
  assign n33 = i0 & i1;
  assign n34 = ~i2 & n33;
  assign n35 = ~i3 & n34;
  assign n36 = ~i4 & n35;
  assign n37 = ~i5 & n36;
  assign n38 = ~i6 & n37;
  assign n39 = i7 & n38;
  assign n40 = i2 & n33;
  assign n41 = i3 & n40;
  assign n42 = ~i4 & n41;
  assign n43 = ~i5 & n42;
  assign n44 = ~i6 & n43;
  assign n45 = ~i7 & n44;
  assign n46 = i3 & n18;
  assign n47 = ~i4 & n46;
  assign n48 = ~i5 & n47;
  assign n49 = ~i6 & n48;
  assign n50 = i7 & n49;
  assign n51 = ~i6 & n28;
  assign n52 = ~i7 & n51;
  assign n53 = i0 & ~i1;
  assign n54 = ~i2 & n53;
  assign n55 = ~i3 & n54;
  assign n56 = ~i4 & n55;
  assign n57 = ~i6 & n56;
  assign n58 = ~i7 & n57;
  assign n59 = ~i3 & n13;
  assign n60 = ~i4 & n59;
  assign n61 = i5 & n60;
  assign n62 = ~i6 & n61;
  assign n63 = ~i7 & n62;
  assign n64 = ~i6 & n46;
  assign n65 = ~i7 & n64;
  assign n66 = ~i0 & i1;
  assign n67 = ~i2 & n66;
  assign n68 = i3 & n67;
  assign n69 = i4 & n68;
  assign n70 = ~i5 & n69;
  assign n71 = ~i6 & n70;
  assign n72 = i7 & n71;
  assign n73 = ~i3 & n67;
  assign n74 = i4 & n73;
  assign n75 = ~i5 & n74;
  assign n76 = ~i6 & n75;
  assign n77 = ~i7 & n76;
  assign n78 = i3 & n54;
  assign n79 = ~i4 & n78;
  assign n80 = i5 & n79;
  assign n81 = ~i6 & n80;
  assign n82 = i7 & n81;
  assign n83 = i4 & n55;
  assign n84 = ~i5 & n83;
  assign n85 = ~i6 & n84;
  assign n86 = ~i7 & n85;
  assign n87 = ~i6 & n35;
  assign n88 = ~i7 & n87;
  assign n89 = i5 & n83;
  assign n90 = ~i6 & n89;
  assign n91 = ~i7 & n90;
  assign n92 = i4 & n78;
  assign n93 = i5 & n92;
  assign n94 = ~i6 & n93;
  assign n95 = i7 & n94;
  assign n96 = ~i5 & n92;
  assign n97 = ~i6 & n96;
  assign n98 = i7 & n97;
  assign n99 = ~i4 & n68;
  assign n100 = ~i6 & n99;
  assign n101 = i7 & n100;
  assign n102 = i5 & n29;
  assign n103 = ~i6 & n102;
  assign n104 = i7 & n103;
  assign n105 = ~n17 & ~n22;
  assign n106 = ~n27 & n105;
  assign n107 = ~n32 & n106;
  assign n108 = ~n39 & n107;
  assign n109 = ~n45 & n108;
  assign n110 = ~n50 & n109;
  assign n111 = ~n52 & n110;
  assign n112 = ~n58 & n111;
  assign n113 = ~n63 & n112;
  assign n114 = ~n65 & n113;
  assign n115 = ~n72 & n114;
  assign n116 = ~n77 & n115;
  assign n117 = ~n82 & n116;
  assign n118 = ~n86 & n117;
  assign n119 = ~n88 & n118;
  assign n120 = ~n91 & n119;
  assign n121 = ~n95 & n120;
  assign n122 = ~n98 & n121;
  assign n123 = ~n101 & n122;
  assign i9 = ~n104 & n123;
  assign n125 = i6 & n13;
  assign n126 = i7 & n125;
  assign n127 = i9 & n126;
  assign n128 = ~i4 & n40;
  assign n129 = ~i5 & n128;
  assign n130 = i6 & n129;
  assign n131 = i7 & n130;
  assign n132 = i9 & n131;
  assign n133 = ~i6 & n13;
  assign n134 = i7 & n133;
  assign n135 = ~i9 & n134;
  assign n136 = ~i6 & n23;
  assign n137 = i7 & n136;
  assign n138 = ~i9 & n137;
  assign n139 = ~i6 & n18;
  assign n140 = i7 & n139;
  assign n141 = ~i9 & n140;
  assign n142 = i4 & n13;
  assign n143 = i6 & n142;
  assign n144 = i7 & n143;
  assign n145 = i9 & n144;
  assign n146 = i4 & n41;
  assign n147 = i6 & n146;
  assign n148 = i7 & n147;
  assign n149 = i9 & n148;
  assign n150 = i4 & n18;
  assign n151 = i6 & n150;
  assign n152 = i7 & n151;
  assign n153 = i9 & n152;
  assign n154 = i4 & n23;
  assign n155 = i6 & n154;
  assign n156 = i7 & n155;
  assign n157 = i9 & n156;
  assign n158 = i1 & i2;
  assign n159 = i3 & n158;
  assign n160 = i4 & n159;
  assign n161 = ~i5 & n160;
  assign n162 = i6 & n161;
  assign n163 = i7 & n162;
  assign n164 = i9 & n163;
  assign n165 = i0 & i2;
  assign n166 = i3 & n165;
  assign n167 = i4 & n166;
  assign n168 = i5 & n167;
  assign n169 = i6 & n168;
  assign n170 = i7 & n169;
  assign n171 = i9 & n170;
  assign n172 = ~i5 & n167;
  assign n173 = i6 & n172;
  assign n174 = i7 & n173;
  assign n175 = i9 & n174;
  assign n176 = ~n70 & ~n145;
  assign n177 = ~n96 & n176;
  assign n178 = ~n93 & n177;
  assign n179 = ~n149 & n178;
  assign n180 = ~n153 & n179;
  assign n181 = ~n157 & n180;
  assign n182 = ~n164 & n181;
  assign n183 = ~n171 & n182;
  assign i10 = ~n175 & n183;
  assign n185 = ~i6 & n142;
  assign n186 = ~i9 & n185;
  assign n187 = i10 & n186;
  assign n188 = i6 & n18;
  assign n189 = i7 & n188;
  assign n190 = i9 & n189;
  assign n191 = ~i5 & n28;
  assign n192 = ~i7 & n191;
  assign n193 = ~i10 & n192;
  assign n194 = ~i6 & n150;
  assign n195 = ~i9 & n194;
  assign n196 = i10 & n195;
  assign n197 = ~i6 & n154;
  assign n198 = ~i9 & n197;
  assign n199 = i10 & n198;
  assign n200 = ~i7 & n92;
  assign n201 = ~i10 & n200;
  assign n202 = i9 & n143;
  assign n203 = i10 & n202;
  assign n204 = i2 & i3;
  assign n205 = ~i4 & n204;
  assign n206 = ~i5 & n205;
  assign n207 = i6 & n206;
  assign n208 = i7 & n207;
  assign n209 = i9 & n208;
  assign n210 = i6 & n23;
  assign n211 = i7 & n210;
  assign n212 = i9 & n211;
  assign n213 = i6 & n41;
  assign n214 = i7 & n213;
  assign n215 = i9 & n214;
  assign n216 = i9 & n151;
  assign n217 = i10 & n216;
  assign n218 = i9 & n155;
  assign n219 = i10 & n218;
  assign n220 = i4 & n158;
  assign n221 = ~i5 & n220;
  assign n222 = i6 & n221;
  assign n223 = ~i7 & n222;
  assign n224 = i9 & n223;
  assign n225 = i10 & n224;
  assign n226 = ~i5 & n204;
  assign n227 = i6 & n226;
  assign n228 = i7 & n227;
  assign n229 = i9 & n228;
  assign n230 = ~i10 & n229;
  assign n231 = i9 & n173;
  assign n232 = i10 & n231;
  assign n233 = i4 & n204;
  assign n234 = i6 & n233;
  assign n235 = ~i7 & n234;
  assign n236 = i9 & n235;
  assign n237 = i10 & n236;
  assign n238 = i4 & n165;
  assign n239 = ~i5 & n238;
  assign n240 = i6 & n239;
  assign n241 = ~i7 & n240;
  assign n242 = i9 & n241;
  assign n243 = i10 & n242;
  assign n244 = i6 & n167;
  assign n245 = i7 & n244;
  assign n246 = i9 & n245;
  assign n247 = ~i10 & n246;
  assign n248 = i4 & n40;
  assign n249 = i6 & n248;
  assign n250 = ~i7 & n249;
  assign n251 = i9 & n250;
  assign n252 = i10 & n251;
  assign n253 = i5 & n238;
  assign n254 = i6 & n253;
  assign n255 = ~i7 & n254;
  assign n256 = i9 & n255;
  assign n257 = i10 & n256;
  assign n258 = i5 & n205;
  assign n259 = i6 & n258;
  assign n260 = i7 & n259;
  assign n261 = i9 & n260;
  assign n262 = i10 & n261;
  assign n263 = ~n127 & ~n132;
  assign n264 = ~n135 & n263;
  assign n265 = ~n138 & n264;
  assign n266 = ~n141 & n265;
  assign n267 = ~n187 & n266;
  assign n268 = ~n190 & n267;
  assign n269 = ~n193 & ~n268;
  assign n270 = ~n135 & ~n269;
  assign n271 = ~n187 & n270;
  assign n272 = ~n141 & n271;
  assign n273 = ~n196 & n272;
  assign n274 = ~n199 & n273;
  assign n275 = ~n201 & ~n274;
  assign n276 = ~n203 & ~n275;
  assign n277 = ~n209 & n276;
  assign n278 = ~n212 & n277;
  assign n279 = ~n196 & n278;
  assign n280 = ~n215 & n279;
  assign n281 = ~n141 & n280;
  assign n282 = ~n141 & n281;
  assign n283 = ~n217 & n282;
  assign n284 = ~n219 & n283;
  assign n285 = ~n135 & n284;
  assign n286 = ~n225 & n285;
  assign n287 = ~n135 & n286;
  assign n288 = ~n230 & n287;
  assign n289 = ~n232 & n288;
  assign n290 = ~n237 & n289;
  assign n291 = ~n243 & n290;
  assign n292 = ~n247 & n291;
  assign n293 = ~n252 & n292;
  assign n294 = ~n257 & n293;
  assign i8 = ~n262 & n294;
  assign n296 = ~i4 & n158;
  assign n297 = i5 & n296;
  assign n298 = i6 & n297;
  assign n299 = ~i7 & n298;
  assign n300 = i8 & n299;
  assign n301 = i9 & n300;
  assign n302 = i10 & n301;
  assign n303 = i5 & n142;
  assign n304 = i6 & n303;
  assign n305 = i7 & n304;
  assign n306 = i9 & n305;
  assign n307 = i5 & n13;
  assign n308 = ~i6 & n307;
  assign n309 = i8 & n308;
  assign n310 = ~i9 & n309;
  assign n311 = i10 & n310;
  assign n312 = i5 & n35;
  assign n313 = ~i7 & n312;
  assign n314 = i8 & n313;
  assign n315 = i10 & n314;
  assign n316 = i6 & n307;
  assign n317 = i8 & n316;
  assign n318 = i9 & n317;
  assign n319 = i10 & n318;
  assign n320 = i4 & n35;
  assign n321 = i5 & n320;
  assign n322 = i7 & n321;
  assign n323 = ~i8 & n322;
  assign n324 = i7 & n316;
  assign n325 = i9 & n324;
  assign n326 = i10 & n325;
  assign n327 = i5 & n99;
  assign n328 = i10 & n327;
  assign n329 = n102 & i10;
  assign n330 = i5 & n146;
  assign n331 = i6 & n330;
  assign n332 = i7 & n331;
  assign n333 = i9 & n332;
  assign n334 = i7 & n312;
  assign n335 = ~i8 & n334;
  assign n336 = i10 & n335;
  assign n337 = i2 & ~i4;
  assign n338 = i5 & n337;
  assign n339 = i6 & n338;
  assign n340 = ~i7 & n339;
  assign n341 = i8 & n340;
  assign n342 = i9 & n341;
  assign n343 = i10 & n342;
  assign n344 = ~i2 & ~i5;
  assign n345 = i2 & ~i5;
  assign n346 = ~i8 & n345;
  assign n347 = ~n344 & ~n346;
  assign n348 = i8 & n345;
  assign n349 = n347 & ~n348;
  assign n350 = ~i1 & i5;
  assign n351 = ~i2 & n350;
  assign n352 = ~i0 & n351;
  assign n353 = i7 & n352;
  assign n354 = n349 & ~n353;
  assign n355 = i0 & n351;
  assign n356 = ~i8 & n355;
  assign n357 = ~i6 & n356;
  assign n358 = ~i3 & n357;
  assign n359 = n354 & ~n358;
  assign n360 = i2 & n350;
  assign n361 = n359 & ~n360;
  assign n362 = i1 & i5;
  assign n363 = n361 & ~n362;
  assign n364 = ~n302 & ~n363;
  assign n365 = ~n306 & n364;
  assign n366 = ~n311 & n365;
  assign n367 = ~n315 & n366;
  assign n368 = ~n319 & n367;
  assign n369 = ~n323 & n368;
  assign n370 = ~n326 & n369;
  assign n371 = ~n328 & n370;
  assign n372 = ~n329 & n371;
  assign n373 = ~n333 & n372;
  assign n374 = ~n336 & n373;
  assign n375 = ~n171 & n374;
  assign n376 = ~n343 & n375;
  assign i11 = ~n262 & n376;
endmodule


