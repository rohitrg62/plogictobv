// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:27:33 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8, i9, i10, i11  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8, i9, i10, i11;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
    n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
    n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
    n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
    n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
    n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
    n97, n98, n99, n100, n102, n103, n104, n105, n106, n107, n108, n109,
    n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
    n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
    n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
    n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
    n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212, n213, n214, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
    n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
    n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n343, n344, n345, n346, n347, n348, n349, n350, n351,
    n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
    n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
    n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
    n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
    n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571;
  assign n13 = i0 & i1;
  assign n14 = i2 & n13;
  assign n15 = i3 & n14;
  assign n16 = i4 & n15;
  assign n17 = i5 & n16;
  assign n18 = i6 & n17;
  assign n19 = i7 & n18;
  assign n20 = ~i2 & n13;
  assign n21 = ~i3 & n20;
  assign n22 = i4 & n21;
  assign n23 = i5 & n22;
  assign n24 = ~i6 & n23;
  assign n25 = i7 & n24;
  assign n26 = ~i0 & i1;
  assign n27 = ~i2 & n26;
  assign n28 = ~i3 & n27;
  assign n29 = i4 & n28;
  assign n30 = ~i5 & n29;
  assign n31 = ~i6 & n30;
  assign n32 = i7 & n31;
  assign n33 = i7 & n30;
  assign n34 = i0 & ~i1;
  assign n35 = ~i2 & n34;
  assign n36 = ~i3 & n35;
  assign n37 = ~i4 & n36;
  assign n38 = ~i5 & n37;
  assign n39 = i6 & n38;
  assign n40 = ~i7 & n39;
  assign n41 = i5 & n37;
  assign n42 = i6 & n41;
  assign n43 = ~i7 & n42;
  assign n44 = i7 & n42;
  assign n45 = ~i4 & n21;
  assign n46 = ~i5 & n45;
  assign n47 = i6 & n46;
  assign n48 = i7 & n47;
  assign n49 = ~i7 & n47;
  assign n50 = i3 & n27;
  assign n51 = i4 & n50;
  assign n52 = ~i5 & n51;
  assign n53 = i6 & n52;
  assign n54 = i7 & n53;
  assign n55 = i3 & n13;
  assign n56 = i4 & n55;
  assign n57 = i5 & n56;
  assign n58 = i6 & n57;
  assign n59 = i7 & n58;
  assign n60 = ~i6 & n41;
  assign n61 = i7 & n60;
  assign n62 = i6 & n23;
  assign n63 = ~i7 & n62;
  assign n64 = ~i0 & ~i1;
  assign n65 = ~i2 & n64;
  assign n66 = i3 & n65;
  assign n67 = i4 & n66;
  assign n68 = ~i5 & n67;
  assign n69 = i6 & n68;
  assign n70 = ~i7 & n69;
  assign n71 = ~i4 & n50;
  assign n72 = i5 & n71;
  assign n73 = i6 & n72;
  assign n74 = i7 & n73;
  assign n75 = i3 & n35;
  assign n76 = ~i4 & n75;
  assign n77 = i5 & n76;
  assign n78 = i6 & n77;
  assign n79 = i7 & n78;
  assign n80 = i5 & n67;
  assign n81 = i6 & n80;
  assign n82 = ~i7 & n81;
  assign n83 = i7 & n81;
  assign n84 = i1 & ~n19;
  assign n85 = ~n25 & n84;
  assign n86 = ~n32 & n85;
  assign n87 = ~n33 & n86;
  assign n88 = ~n40 & ~n87;
  assign n89 = ~n43 & n88;
  assign n90 = ~n44 & n89;
  assign n91 = ~n48 & ~n90;
  assign n92 = ~n49 & n91;
  assign n93 = ~n54 & n92;
  assign n94 = ~n59 & n93;
  assign n95 = ~n61 & ~n94;
  assign n96 = ~n63 & ~n95;
  assign n97 = ~n70 & ~n96;
  assign n98 = ~n74 & ~n97;
  assign n99 = ~n79 & ~n98;
  assign n100 = ~n82 & n99;
  assign i10 = n83 | ~n100;
  assign n102 = i4 & n36;
  assign n103 = i5 & n102;
  assign n104 = i6 & n103;
  assign n105 = i7 & n104;
  assign n106 = ~i10 & n105;
  assign n107 = ~i3 & n65;
  assign n108 = i4 & n107;
  assign n109 = ~i5 & n108;
  assign n110 = ~i6 & n109;
  assign n111 = ~i10 & n110;
  assign n112 = i1 & ~i2;
  assign n113 = ~i3 & n112;
  assign n114 = i4 & n113;
  assign n115 = i5 & n114;
  assign n116 = ~i6 & n115;
  assign n117 = i7 & n116;
  assign n118 = ~i10 & n117;
  assign n119 = n32 & ~i10;
  assign n120 = ~i3 & n14;
  assign n121 = i4 & n120;
  assign n122 = i5 & n121;
  assign n123 = i6 & n122;
  assign n124 = ~i7 & n123;
  assign n125 = i10 & n124;
  assign n126 = i6 & n30;
  assign n127 = i7 & n126;
  assign n128 = ~i10 & n127;
  assign n129 = ~i0 & ~i2;
  assign n130 = ~i3 & n129;
  assign n131 = i4 & n130;
  assign n132 = i5 & n131;
  assign n133 = ~i6 & n132;
  assign n134 = ~i10 & n133;
  assign n135 = n62 & i10;
  assign n136 = i5 & n45;
  assign n137 = i6 & n136;
  assign n138 = ~i7 & n137;
  assign n139 = i10 & n138;
  assign n140 = i2 & n34;
  assign n141 = i3 & n140;
  assign n142 = i4 & n141;
  assign n143 = ~i5 & n142;
  assign n144 = i6 & n143;
  assign n145 = i7 & n144;
  assign n146 = ~i10 & n145;
  assign n147 = ~i7 & n126;
  assign n148 = i10 & n147;
  assign n149 = n43 & i10;
  assign n150 = n54 & ~i10;
  assign n151 = i5 & n51;
  assign n152 = i6 & n151;
  assign n153 = ~i7 & n152;
  assign n154 = i10 & n153;
  assign n155 = n49 & ~i10;
  assign n156 = n61 & i10;
  assign n157 = i2 & n26;
  assign n158 = i3 & n157;
  assign n159 = ~i4 & n158;
  assign n160 = i5 & n159;
  assign n161 = i6 & n160;
  assign n162 = i7 & n161;
  assign n163 = i10 & n162;
  assign n164 = i7 & n39;
  assign n165 = ~i10 & n164;
  assign n166 = n70 & i10;
  assign n167 = i7 & n69;
  assign n168 = ~i10 & n167;
  assign n169 = ~i4 & n66;
  assign n170 = i5 & n169;
  assign n171 = i6 & n170;
  assign n172 = ~i7 & n171;
  assign n173 = ~i10 & n172;
  assign n174 = n79 & i10;
  assign n175 = ~i5 & n102;
  assign n176 = i6 & n175;
  assign n177 = i7 & n176;
  assign n178 = ~i10 & n177;
  assign n179 = n82 & i10;
  assign n180 = ~i6 & i7;
  assign n181 = ~i10 & n180;
  assign n182 = ~i5 & i6;
  assign n183 = ~i2 & n182;
  assign n184 = i10 & n183;
  assign n185 = ~i3 & n184;
  assign n186 = ~i7 & n185;
  assign n187 = ~n181 & ~n186;
  assign n188 = i3 & n184;
  assign n189 = n187 & ~n188;
  assign n190 = i2 & n182;
  assign n191 = n189 & ~n190;
  assign n192 = ~n106 & n191;
  assign n193 = ~n111 & ~n192;
  assign n194 = ~n118 & ~n193;
  assign n195 = ~n119 & n194;
  assign n196 = ~n125 & n195;
  assign n197 = ~n128 & n196;
  assign n198 = ~n134 & ~n197;
  assign n199 = ~n135 & ~n198;
  assign n200 = ~n139 & n199;
  assign n201 = ~n146 & ~n200;
  assign n202 = ~n148 & n201;
  assign n203 = ~n149 & ~n202;
  assign n204 = ~n150 & ~n203;
  assign n205 = ~n154 & ~n204;
  assign n206 = ~n155 & n205;
  assign n207 = ~n156 & ~n206;
  assign n208 = ~n163 & ~n207;
  assign n209 = ~n165 & n208;
  assign n210 = ~n166 & n209;
  assign n211 = ~n168 & n210;
  assign n212 = ~n173 & n211;
  assign n213 = ~n174 & n212;
  assign n214 = ~n178 & n213;
  assign i11 = n179 | ~n214;
  assign n216 = ~i4 & n130;
  assign n217 = i5 & n216;
  assign n218 = ~i6 & n217;
  assign n219 = i7 & n218;
  assign n220 = i10 & n219;
  assign n221 = ~i4 & n28;
  assign n222 = i5 & n221;
  assign n223 = i6 & n222;
  assign n224 = ~i7 & n223;
  assign n225 = i10 & n224;
  assign n226 = ~i11 & n225;
  assign n227 = i7 & n137;
  assign n228 = i10 & n227;
  assign n229 = ~i11 & n228;
  assign n230 = n19 & ~i10;
  assign n231 = ~i11 & n230;
  assign n232 = ~i4 & n107;
  assign n233 = ~i5 & n232;
  assign n234 = ~i6 & n233;
  assign n235 = i7 & n234;
  assign n236 = ~i10 & n235;
  assign n237 = i11 & n236;
  assign n238 = n118 & i11;
  assign n239 = i5 & n29;
  assign n240 = ~i6 & n239;
  assign n241 = ~i7 & n240;
  assign n242 = i10 & n241;
  assign n243 = ~i1 & ~i2;
  assign n244 = ~i3 & n243;
  assign n245 = i4 & n244;
  assign n246 = ~i5 & n245;
  assign n247 = ~i6 & n246;
  assign n248 = i7 & n247;
  assign n249 = ~i10 & n248;
  assign n250 = i11 & n249;
  assign n251 = i7 & n23;
  assign n252 = i10 & n251;
  assign n253 = i11 & n252;
  assign n254 = i6 & n239;
  assign n255 = i10 & n254;
  assign n256 = ~i11 & n255;
  assign n257 = i5 & n107;
  assign n258 = n139 & i11;
  assign n259 = n145 & ~i11;
  assign n260 = i7 & n152;
  assign n261 = i10 & n260;
  assign n262 = ~i11 & n261;
  assign n263 = n154 & i11;
  assign n264 = i0 & ~i2;
  assign n265 = ~i3 & n264;
  assign n266 = ~i4 & n265;
  assign n267 = ~i5 & n266;
  assign n268 = i6 & n267;
  assign n269 = ~i7 & n268;
  assign n270 = i10 & n269;
  assign n271 = i11 & n270;
  assign n272 = n59 & ~i10;
  assign n273 = ~i11 & n272;
  assign n274 = ~i10 & n176;
  assign n275 = ~i11 & n274;
  assign n276 = n62 & ~i10;
  assign n277 = i11 & n276;
  assign n278 = n166 & i11;
  assign n279 = i5 & n50;
  assign n280 = i6 & n279;
  assign n281 = i7 & n280;
  assign n282 = ~i10 & n281;
  assign n283 = ~i11 & n282;
  assign n284 = ~i5 & n66;
  assign n285 = i6 & n284;
  assign n286 = i7 & n285;
  assign n287 = ~i11 & n286;
  assign n288 = i4 & n75;
  assign n289 = ~i5 & n288;
  assign n290 = i6 & n289;
  assign n291 = i7 & n290;
  assign n292 = ~i10 & n291;
  assign n293 = ~i11 & n292;
  assign n294 = i7 & n175;
  assign n295 = ~i10 & n294;
  assign n296 = i11 & n295;
  assign n297 = ~i10 & ~i11;
  assign n298 = ~i4 & n297;
  assign n299 = i6 & n298;
  assign n300 = i4 & n297;
  assign n301 = ~i0 & n300;
  assign n302 = ~i3 & n301;
  assign n303 = ~n299 & ~n302;
  assign n304 = i3 & n301;
  assign n305 = ~i6 & n304;
  assign n306 = ~i7 & n305;
  assign n307 = n303 & ~n306;
  assign n308 = i6 & n304;
  assign n309 = n307 & ~n308;
  assign n310 = i0 & n300;
  assign n311 = ~i6 & n310;
  assign n312 = n309 & ~n311;
  assign n313 = i6 & n310;
  assign n314 = ~i1 & n313;
  assign n315 = n312 & ~n314;
  assign n316 = ~i10 & i11;
  assign n317 = n315 & ~n316;
  assign n318 = ~i10 & n317;
  assign n319 = ~n220 & ~n318;
  assign n320 = ~n226 & n319;
  assign n321 = ~n229 & n320;
  assign n322 = ~n231 & n321;
  assign n323 = ~n237 & n322;
  assign n324 = ~n238 & n323;
  assign n325 = ~n242 & n324;
  assign n326 = ~n250 & n325;
  assign n327 = ~n253 & n326;
  assign n328 = ~n256 & n327;
  assign n329 = ~n257 & ~n328;
  assign n330 = ~n258 & ~n329;
  assign n331 = ~n259 & n330;
  assign n332 = ~n262 & n331;
  assign n333 = ~n263 & n332;
  assign n334 = ~n271 & n333;
  assign n335 = ~n273 & n334;
  assign n336 = ~n275 & n335;
  assign n337 = ~n277 & n336;
  assign n338 = ~n278 & n337;
  assign n339 = ~n283 & n338;
  assign n340 = ~n287 & n339;
  assign n341 = ~n293 & n340;
  assign i9 = ~n296 & n341;
  assign n343 = ~i4 & n27;
  assign n344 = i5 & n343;
  assign n345 = ~i6 & n344;
  assign n346 = i7 & n345;
  assign n347 = i9 & n346;
  assign n348 = i10 & n347;
  assign n349 = ~i11 & n348;
  assign n350 = i5 & n130;
  assign n351 = ~i6 & n350;
  assign n352 = i7 & n351;
  assign n353 = i10 & n352;
  assign n354 = i6 & n217;
  assign n355 = ~i7 & n354;
  assign n356 = ~i9 & n355;
  assign n357 = i10 & n356;
  assign n358 = ~i5 & n22;
  assign n359 = i6 & n358;
  assign n360 = i7 & n359;
  assign n361 = i9 & n360;
  assign n362 = i10 & n361;
  assign n363 = ~i11 & n362;
  assign n364 = n105 & i9;
  assign n365 = ~i10 & n364;
  assign n366 = i11 & n365;
  assign n367 = n227 & ~i9;
  assign n368 = i10 & n367;
  assign n369 = ~i11 & n368;
  assign n370 = i4 & n20;
  assign n371 = i5 & n370;
  assign n372 = ~i6 & n371;
  assign n373 = i7 & n372;
  assign n374 = i9 & n373;
  assign n375 = i10 & n374;
  assign n376 = ~i11 & n375;
  assign n377 = ~i7 & n116;
  assign n378 = i9 & n377;
  assign n379 = i10 & n378;
  assign n380 = ~i11 & n379;
  assign n381 = ~i3 & n13;
  assign n382 = i4 & n381;
  assign n383 = i5 & n382;
  assign n384 = i6 & n383;
  assign n385 = ~i7 & n384;
  assign n386 = i9 & n385;
  assign n387 = i10 & n386;
  assign n388 = i11 & n387;
  assign n389 = n127 & i9;
  assign n390 = ~i10 & n389;
  assign n391 = i11 & n390;
  assign n392 = n133 & ~i9;
  assign n393 = i10 & n392;
  assign n394 = n175 & i9;
  assign n395 = ~i10 & n394;
  assign n396 = ~i11 & n395;
  assign n397 = ~i5 & n221;
  assign n398 = i6 & n397;
  assign n399 = i7 & n398;
  assign n400 = i9 & n399;
  assign n401 = i10 & n400;
  assign n402 = ~i11 & n401;
  assign n403 = ~i2 & ~i3;
  assign n404 = ~i4 & n403;
  assign n405 = ~i5 & n404;
  assign n406 = i6 & n405;
  assign n407 = ~i7 & n406;
  assign n408 = i9 & n407;
  assign n409 = i10 & n408;
  assign n410 = i11 & n409;
  assign n411 = n145 & ~i9;
  assign n412 = ~i10 & n411;
  assign n413 = ~i11 & n412;
  assign n414 = i3 & n129;
  assign n415 = i4 & n414;
  assign n416 = i5 & n415;
  assign n417 = i6 & n416;
  assign n418 = i7 & n417;
  assign n419 = ~i9 & n418;
  assign n420 = i10 & n419;
  assign n421 = ~i11 & n420;
  assign n422 = n147 & i9;
  assign n423 = i10 & n422;
  assign n424 = n44 & i9;
  assign n425 = i10 & n424;
  assign n426 = ~i11 & n425;
  assign n427 = n48 & i9;
  assign n428 = ~i10 & n427;
  assign n429 = ~i11 & n428;
  assign n430 = n54 & i9;
  assign n431 = ~i10 & n430;
  assign n432 = ~i11 & n431;
  assign n433 = ~i2 & i3;
  assign n434 = i4 & n433;
  assign n435 = i5 & n434;
  assign n436 = i6 & n435;
  assign n437 = i7 & n436;
  assign n438 = ~i9 & n437;
  assign n439 = ~i10 & n438;
  assign n440 = ~i11 & n439;
  assign n441 = ~i3 & n140;
  assign n442 = i4 & n441;
  assign n443 = ~i5 & n442;
  assign n444 = i6 & n443;
  assign n445 = ~i7 & n444;
  assign n446 = i9 & n445;
  assign n447 = ~i10 & n446;
  assign n448 = i11 & n447;
  assign n449 = i4 & n265;
  assign n450 = i5 & n449;
  assign n451 = i6 & n450;
  assign n452 = ~i7 & n451;
  assign n453 = i9 & n452;
  assign n454 = ~i10 & n453;
  assign n455 = ~i11 & n454;
  assign n456 = i3 & n26;
  assign n457 = ~i4 & n456;
  assign n458 = i5 & n457;
  assign n459 = i6 & n458;
  assign n460 = i7 & n459;
  assign n461 = i9 & n460;
  assign n462 = i10 & n461;
  assign n463 = i11 & n462;
  assign n464 = i6 & n115;
  assign n465 = ~i7 & n464;
  assign n466 = ~i10 & n465;
  assign n467 = i11 & n466;
  assign n468 = i6 & n67;
  assign n469 = ~i7 & n468;
  assign n470 = i10 & n469;
  assign n471 = i11 & n470;
  assign n472 = n167 & i9;
  assign n473 = ~i10 & n472;
  assign n474 = i11 & n473;
  assign n475 = i5 & n414;
  assign n476 = i6 & n475;
  assign n477 = i7 & n476;
  assign n478 = ~i9 & n477;
  assign n479 = ~i10 & n478;
  assign n480 = ~i11 & n479;
  assign n481 = n172 & i9;
  assign n482 = ~i10 & n481;
  assign n483 = i11 & n482;
  assign n484 = i3 & n243;
  assign n485 = ~i4 & n484;
  assign n486 = i5 & n485;
  assign n487 = i6 & n486;
  assign n488 = i7 & n487;
  assign n489 = i9 & n488;
  assign n490 = i10 & n489;
  assign n491 = i11 & n490;
  assign n492 = i6 & n246;
  assign n493 = ~i9 & n492;
  assign n494 = ~i10 & n493;
  assign n495 = ~i11 & n494;
  assign n496 = i9 & n469;
  assign n497 = i10 & n496;
  assign n498 = i11 & n497;
  assign n499 = i9 & n418;
  assign n500 = i10 & n499;
  assign n501 = ~i11 & n500;
  assign n502 = ~i9 & n464;
  assign n503 = ~i10 & n502;
  assign n504 = ~i11 & n503;
  assign n505 = i4 & n484;
  assign n506 = i6 & n505;
  assign n507 = i7 & n506;
  assign n508 = ~i9 & n507;
  assign n509 = ~i10 & n508;
  assign n510 = ~i11 & n509;
  assign n511 = i6 & n414;
  assign n512 = i7 & n511;
  assign n513 = ~i9 & n512;
  assign n514 = ~i10 & n513;
  assign n515 = ~i11 & n514;
  assign n516 = ~i6 & ~i9;
  assign n517 = i11 & n516;
  assign n518 = i10 & n517;
  assign n519 = ~i3 & i9;
  assign n520 = ~i0 & n519;
  assign n521 = ~i7 & n520;
  assign n522 = ~i1 & n521;
  assign n523 = i11 & n522;
  assign n524 = ~n518 & ~n523;
  assign n525 = i1 & n521;
  assign n526 = ~i6 & n525;
  assign n527 = n524 & ~n526;
  assign n528 = i6 & n525;
  assign n529 = n527 & ~n528;
  assign n530 = i3 & i9;
  assign n531 = ~i10 & n530;
  assign n532 = n529 & ~n531;
  assign n533 = i10 & n530;
  assign n534 = ~i1 & n533;
  assign n535 = ~i5 & n534;
  assign n536 = n532 & ~n535;
  assign n537 = ~n349 & n536;
  assign n538 = ~n353 & ~n537;
  assign n539 = ~n357 & n538;
  assign n540 = ~n363 & ~n539;
  assign n541 = ~n366 & n540;
  assign n542 = ~n369 & n541;
  assign n543 = ~n376 & n542;
  assign n544 = ~n380 & n543;
  assign n545 = ~n388 & n544;
  assign n546 = ~n391 & n545;
  assign n547 = ~n393 & ~n546;
  assign n548 = ~n396 & ~n547;
  assign n549 = ~n402 & n548;
  assign n550 = ~n410 & ~n549;
  assign n551 = ~n413 & n550;
  assign n552 = ~n421 & ~n551;
  assign n553 = ~n423 & ~n552;
  assign n554 = ~n426 & ~n553;
  assign n555 = ~n429 & n554;
  assign n556 = ~n432 & n555;
  assign n557 = ~n440 & n556;
  assign n558 = ~n448 & n557;
  assign n559 = ~n455 & n558;
  assign n560 = ~n463 & n559;
  assign n561 = ~n467 & ~n560;
  assign n562 = ~n471 & n561;
  assign n563 = ~n474 & n562;
  assign n564 = ~n480 & ~n563;
  assign n565 = ~n483 & ~n564;
  assign n566 = ~n491 & n565;
  assign n567 = ~n495 & ~n566;
  assign n568 = ~n498 & ~n567;
  assign n569 = ~n501 & ~n568;
  assign n570 = ~n504 & n569;
  assign n571 = ~n510 & n570;
  assign i8 = n515 | ~n571;
endmodule


