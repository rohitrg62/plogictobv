// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 15:53:31 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8;
  assign i8 = 1'b1;
endmodule


