// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:26:54 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8, i9, i10, i11  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8, i9, i10, i11;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
    n27, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
    n42, n43, n44, n45, n46, n47, n48, n49, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
    n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306;
  assign n13 = i0 & i1;
  assign n14 = i2 & n13;
  assign n15 = i3 & n14;
  assign n16 = i4 & n15;
  assign n17 = i5 & n16;
  assign n18 = ~i6 & n17;
  assign n19 = i7 & n18;
  assign n20 = ~i6 & n16;
  assign n21 = i7 & n20;
  assign n22 = ~i0 & i2;
  assign n23 = i2 & ~n22;
  assign n24 = i0 & i2;
  assign n25 = ~i6 & n24;
  assign n26 = n23 & ~n25;
  assign n27 = ~n19 & ~n26;
  assign i11 = ~n21 & n27;
  assign n29 = n19 & ~i11;
  assign n30 = i5 & n15;
  assign n31 = ~i6 & n30;
  assign n32 = i7 & n31;
  assign n33 = i11 & n32;
  assign n34 = ~i6 & n15;
  assign n35 = i7 & n34;
  assign n36 = i11 & n35;
  assign n37 = ~i3 & ~i11;
  assign n38 = ~i1 & n37;
  assign n39 = ~i3 & i11;
  assign n40 = ~i7 & n39;
  assign n41 = ~n38 & ~n40;
  assign n42 = i3 & i11;
  assign n43 = ~i0 & n42;
  assign n44 = n41 & ~n43;
  assign n45 = i0 & n42;
  assign n46 = i2 & n45;
  assign n47 = n44 & ~n46;
  assign n48 = ~n29 & ~n47;
  assign n49 = ~n33 & n48;
  assign i10 = ~n36 & n49;
  assign n51 = ~i0 & ~i1;
  assign n52 = i2 & n51;
  assign n53 = i3 & n52;
  assign n54 = i6 & n53;
  assign n55 = ~i7 & n54;
  assign n56 = i10 & n55;
  assign n57 = i11 & n56;
  assign n58 = i0 & ~i1;
  assign n59 = ~i2 & n58;
  assign n60 = i3 & n59;
  assign n61 = ~i4 & n60;
  assign n62 = ~i6 & n61;
  assign n63 = i7 & n62;
  assign n64 = ~i10 & n63;
  assign n65 = i11 & n64;
  assign n66 = ~i2 & n13;
  assign n67 = i3 & n66;
  assign n68 = ~i5 & n67;
  assign n69 = ~i6 & n68;
  assign n70 = i7 & n69;
  assign n71 = ~i10 & n70;
  assign n72 = i11 & n71;
  assign n73 = ~i0 & i1;
  assign n74 = i2 & n73;
  assign n75 = ~i3 & n74;
  assign n76 = ~i6 & n75;
  assign n77 = i7 & n76;
  assign n78 = ~i10 & n77;
  assign n79 = i11 & n78;
  assign n80 = i4 & n75;
  assign n81 = i5 & n80;
  assign n82 = ~i6 & n81;
  assign n83 = i10 & n82;
  assign n84 = i11 & n83;
  assign n85 = ~i3 & n52;
  assign n86 = i5 & n85;
  assign n87 = ~i6 & n86;
  assign n88 = i7 & n87;
  assign n89 = ~i10 & n88;
  assign n90 = i11 & n89;
  assign n91 = ~i4 & n75;
  assign n92 = ~i5 & n91;
  assign n93 = i6 & n92;
  assign n94 = ~i7 & n93;
  assign n95 = i10 & n94;
  assign n96 = i11 & n95;
  assign n97 = ~i4 & n67;
  assign n98 = i5 & n97;
  assign n99 = ~i6 & n98;
  assign n100 = i7 & n99;
  assign n101 = ~i10 & n100;
  assign n102 = i11 & n101;
  assign n103 = i4 & n67;
  assign n104 = ~i6 & n103;
  assign n105 = ~i7 & n104;
  assign n106 = ~i10 & n105;
  assign n107 = i11 & n106;
  assign n108 = ~i6 & n85;
  assign n109 = i7 & n108;
  assign n110 = ~i10 & n109;
  assign n111 = i11 & n110;
  assign n112 = i4 & n60;
  assign n113 = i5 & n112;
  assign n114 = ~i6 & n113;
  assign n115 = ~i7 & n114;
  assign n116 = ~i10 & n115;
  assign n117 = i11 & n116;
  assign n118 = i5 & n60;
  assign n119 = ~i6 & n118;
  assign n120 = ~i7 & n119;
  assign n121 = ~i10 & n120;
  assign n122 = i11 & n121;
  assign n123 = i4 & n85;
  assign n124 = ~i6 & n123;
  assign n125 = i10 & n124;
  assign n126 = i11 & n125;
  assign n127 = i4 & n52;
  assign n128 = i5 & n127;
  assign n129 = ~i6 & n128;
  assign n130 = i7 & n129;
  assign n131 = i10 & n130;
  assign n132 = i11 & n131;
  assign n133 = ~i6 & n112;
  assign n134 = ~i7 & n133;
  assign n135 = ~i10 & n134;
  assign n136 = i11 & n135;
  assign n137 = ~i6 & n80;
  assign n138 = i10 & n137;
  assign n139 = i11 & n138;
  assign n140 = i3 & n22;
  assign n141 = i6 & n140;
  assign n142 = ~i7 & n141;
  assign n143 = i10 & n142;
  assign n144 = i11 & n143;
  assign n145 = ~i3 & n24;
  assign n146 = ~i4 & n145;
  assign n147 = i6 & n146;
  assign n148 = ~i7 & n147;
  assign n149 = i10 & n148;
  assign n150 = ~i11 & n149;
  assign n151 = i5 & n53;
  assign n152 = ~i6 & n151;
  assign n153 = i7 & n152;
  assign n154 = i10 & n153;
  assign n155 = i11 & n154;
  assign n156 = i3 & n74;
  assign n157 = ~i4 & n156;
  assign n158 = ~i5 & n157;
  assign n159 = i6 & n158;
  assign n160 = i10 & n159;
  assign n161 = i11 & n160;
  assign n162 = i4 & n156;
  assign n163 = ~i6 & n162;
  assign n164 = i7 & n163;
  assign n165 = i10 & n164;
  assign n166 = i11 & n165;
  assign n167 = i4 & n53;
  assign n168 = ~i6 & n167;
  assign n169 = i7 & n168;
  assign n170 = i10 & n169;
  assign n171 = i11 & n170;
  assign n172 = i1 & i2;
  assign n173 = i3 & n172;
  assign n174 = i4 & n173;
  assign n175 = i5 & n174;
  assign n176 = ~i6 & n175;
  assign n177 = i7 & n176;
  assign n178 = ~i10 & n177;
  assign n179 = ~i11 & n178;
  assign n180 = ~i11 & ~i10;
  assign n181 = ~i2 & n180;
  assign n182 = i5 & n181;
  assign n183 = i6 & n182;
  assign n184 = ~i11 & i10;
  assign n185 = ~i6 & n184;
  assign n186 = ~n183 & ~n185;
  assign n187 = i0 & i11;
  assign n188 = ~i2 & n187;
  assign n189 = i10 & n188;
  assign n190 = n186 & ~n189;
  assign n191 = i2 & n187;
  assign n192 = n190 & ~n191;
  assign n193 = ~n57 & n192;
  assign n194 = ~n65 & n193;
  assign n195 = ~n72 & n194;
  assign n196 = ~n79 & n195;
  assign n197 = ~n84 & n196;
  assign n198 = ~n90 & n197;
  assign n199 = ~n96 & n198;
  assign n200 = ~n102 & n199;
  assign n201 = ~n107 & n200;
  assign n202 = ~n111 & n201;
  assign n203 = ~n117 & n202;
  assign n204 = ~n122 & n203;
  assign n205 = ~n126 & n204;
  assign n206 = ~n132 & n205;
  assign n207 = ~n136 & n206;
  assign n208 = ~n139 & n207;
  assign n209 = ~n144 & n208;
  assign n210 = ~n150 & n209;
  assign n211 = ~n155 & n210;
  assign n212 = ~n161 & n211;
  assign n213 = ~n166 & n212;
  assign n214 = ~n171 & n213;
  assign i9 = ~n179 & ~n214;
  assign n216 = ~i2 & n51;
  assign n217 = i3 & n216;
  assign n218 = i4 & n217;
  assign n219 = ~i6 & n218;
  assign n220 = ~i7 & n219;
  assign n221 = ~i9 & n220;
  assign n222 = i10 & n221;
  assign n223 = i11 & n222;
  assign n224 = ~i2 & n73;
  assign n225 = i3 & n224;
  assign n226 = ~i4 & n225;
  assign n227 = ~i5 & n226;
  assign n228 = ~i6 & n227;
  assign n229 = i7 & n228;
  assign n230 = ~i9 & n229;
  assign n231 = i10 & n230;
  assign n232 = i11 & n231;
  assign n233 = ~i6 & n67;
  assign n234 = ~i7 & n233;
  assign n235 = ~i9 & n234;
  assign n236 = ~i10 & n235;
  assign n237 = i11 & n236;
  assign n238 = i4 & n225;
  assign n239 = ~i6 & n238;
  assign n240 = ~i7 & n239;
  assign n241 = ~i9 & n240;
  assign n242 = i10 & n241;
  assign n243 = i11 & n242;
  assign n244 = i2 & i3;
  assign n245 = i6 & n244;
  assign n246 = ~i7 & n245;
  assign n247 = i9 & n246;
  assign n248 = ~i4 & n173;
  assign n249 = ~i5 & n248;
  assign n250 = i6 & n249;
  assign n251 = i9 & n250;
  assign n252 = n18 & i9;
  assign n253 = n87 & ~i9;
  assign n254 = i10 & n253;
  assign n255 = i11 & n254;
  assign n256 = ~i6 & n173;
  assign n257 = i7 & n256;
  assign n258 = i9 & n257;
  assign n259 = ~i10 & n258;
  assign n260 = n20 & i9;
  assign n261 = i11 & n260;
  assign n262 = n31 & i9;
  assign n263 = i10 & n262;
  assign n264 = n34 & i9;
  assign n265 = i10 & n264;
  assign n266 = i11 & n265;
  assign n267 = ~i10 & ~i9;
  assign n268 = i11 & n267;
  assign n269 = ~i1 & n268;
  assign n270 = ~i6 & n269;
  assign n271 = i6 & n269;
  assign n272 = ~n270 & ~n271;
  assign n273 = i1 & n268;
  assign n274 = i2 & n273;
  assign n275 = n272 & ~n274;
  assign n276 = i10 & ~i9;
  assign n277 = ~i6 & n276;
  assign n278 = ~i2 & n277;
  assign n279 = i5 & n278;
  assign n280 = n275 & ~n279;
  assign n281 = i2 & n277;
  assign n282 = n280 & ~n281;
  assign n283 = i6 & n276;
  assign n284 = ~i11 & n283;
  assign n285 = ~i1 & n284;
  assign n286 = n282 & ~n285;
  assign n287 = i1 & n284;
  assign n288 = n286 & ~n287;
  assign n289 = i11 & n283;
  assign n290 = ~i5 & n289;
  assign n291 = ~i4 & n290;
  assign n292 = ~i1 & n291;
  assign n293 = n288 & ~n292;
  assign n294 = ~i9 & n293;
  assign n295 = ~n223 & n294;
  assign n296 = ~n232 & n295;
  assign n297 = ~n237 & n296;
  assign n298 = ~n243 & n297;
  assign n299 = ~n247 & n298;
  assign n300 = ~n251 & n299;
  assign n301 = ~n252 & ~n300;
  assign n302 = ~n255 & n301;
  assign n303 = ~n259 & n302;
  assign n304 = ~n259 & n303;
  assign n305 = ~n261 & n304;
  assign n306 = ~n263 & n305;
  assign i8 = ~n266 & n306;
endmodule


