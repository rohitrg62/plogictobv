// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:27:57 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8, i9, i10, i11  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8, i9, i10, i11;
  wire n13, n14, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
    n28, n29, n30, n31, n32, n33, n35, n36, n37, n38, n39, n40, n41, n42,
    n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
    n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320;
  assign n13 = ~i1 & ~i5;
  assign n14 = i1 & i5;
  assign i8 = ~n13 & ~n14;
  assign n16 = i0 & i1;
  assign n17 = ~i4 & n16;
  assign n18 = i8 & n17;
  assign n19 = ~i0 & i1;
  assign n20 = i4 & n19;
  assign n21 = i8 & n20;
  assign n22 = ~i0 & ~i1;
  assign n23 = ~i4 & n22;
  assign n24 = ~i0 & ~i4;
  assign n25 = ~i8 & n24;
  assign n26 = i0 & ~i1;
  assign n27 = i4 & n26;
  assign n28 = i0 & i4;
  assign n29 = ~i8 & n28;
  assign n30 = ~n18 & ~n21;
  assign n31 = ~n23 & n30;
  assign n32 = ~n25 & n31;
  assign n33 = ~n27 & n32;
  assign i9 = ~n29 & n33;
  assign n35 = i2 & n16;
  assign n36 = i3 & n35;
  assign n37 = ~i6 & n36;
  assign n38 = i8 & n37;
  assign n39 = i0 & i2;
  assign n40 = i3 & n39;
  assign n41 = ~i6 & n40;
  assign n42 = i9 & n41;
  assign n43 = i0 & ~i2;
  assign n44 = i3 & n43;
  assign n45 = i6 & n44;
  assign n46 = i9 & n45;
  assign n47 = ~i3 & n39;
  assign n48 = ~i6 & n47;
  assign n49 = ~i7 & n48;
  assign n50 = i9 & n49;
  assign n51 = ~i3 & n43;
  assign n52 = i6 & n51;
  assign n53 = ~i7 & n52;
  assign n54 = i9 & n53;
  assign n55 = i1 & ~i2;
  assign n56 = i3 & n55;
  assign n57 = i6 & n56;
  assign n58 = i8 & n57;
  assign n59 = i9 & n58;
  assign n60 = ~i3 & n55;
  assign n61 = ~i6 & n60;
  assign n62 = i7 & n61;
  assign n63 = i8 & n62;
  assign n64 = i9 & n63;
  assign n65 = i6 & n60;
  assign n66 = ~i7 & n65;
  assign n67 = i8 & n66;
  assign n68 = i9 & n67;
  assign n69 = ~i0 & ~i2;
  assign n70 = i3 & n69;
  assign n71 = ~i6 & n70;
  assign n72 = i7 & n71;
  assign n73 = ~i8 & n72;
  assign n74 = ~i9 & n72;
  assign n75 = ~i3 & n69;
  assign n76 = ~i6 & n75;
  assign n77 = ~i9 & n76;
  assign n78 = ~i2 & n22;
  assign n79 = ~i3 & n78;
  assign n80 = ~i6 & n79;
  assign n81 = i6 & n70;
  assign n82 = ~i7 & n81;
  assign n83 = ~i8 & n82;
  assign n84 = ~i8 & n76;
  assign n85 = i1 & i2;
  assign n86 = i3 & n85;
  assign n87 = ~i6 & n86;
  assign n88 = i8 & n87;
  assign n89 = i9 & n88;
  assign n90 = ~i3 & n85;
  assign n91 = ~i6 & n90;
  assign n92 = ~i7 & n91;
  assign n93 = i8 & n92;
  assign n94 = i9 & n93;
  assign n95 = i2 & n22;
  assign n96 = i3 & n95;
  assign n97 = ~i6 & n96;
  assign n98 = ~i7 & n97;
  assign n99 = i6 & n96;
  assign n100 = i7 & n99;
  assign n101 = ~i3 & n95;
  assign n102 = i6 & n101;
  assign n103 = ~i0 & i2;
  assign n104 = i3 & n103;
  assign n105 = i6 & n104;
  assign n106 = i7 & n105;
  assign n107 = ~i8 & n106;
  assign n108 = ~i3 & n103;
  assign n109 = i6 & n108;
  assign n110 = ~i9 & n109;
  assign n111 = ~i8 & n109;
  assign n112 = i6 & n90;
  assign n113 = i7 & n112;
  assign n114 = i8 & n113;
  assign n115 = i9 & n114;
  assign n116 = ~i1 & ~i2;
  assign n117 = ~i3 & n116;
  assign n118 = ~i6 & n117;
  assign n119 = ~i9 & n118;
  assign n120 = ~i2 & ~i3;
  assign n121 = ~i6 & n120;
  assign n122 = ~i8 & n121;
  assign n123 = ~i9 & n122;
  assign n124 = ~i6 & n51;
  assign n125 = i7 & n124;
  assign n126 = i9 & n125;
  assign n127 = i6 & n47;
  assign n128 = i7 & n127;
  assign n129 = i9 & n128;
  assign n130 = ~i2 & n16;
  assign n131 = ~i3 & n130;
  assign n132 = i6 & n131;
  assign n133 = ~i7 & n132;
  assign n134 = i8 & n133;
  assign n135 = i3 & n116;
  assign n136 = i6 & n135;
  assign n137 = ~i7 & n136;
  assign n138 = ~i9 & n137;
  assign n139 = ~i6 & n131;
  assign n140 = i7 & n139;
  assign n141 = i8 & n140;
  assign n142 = ~i3 & n35;
  assign n143 = ~i6 & n142;
  assign n144 = ~i7 & n143;
  assign n145 = i8 & n144;
  assign n146 = ~i1 & i2;
  assign n147 = ~i3 & n146;
  assign n148 = i6 & n147;
  assign n149 = ~i9 & n148;
  assign n150 = i6 & n142;
  assign n151 = i7 & n150;
  assign n152 = i8 & n151;
  assign n153 = ~i9 & n106;
  assign n154 = i3 & n78;
  assign n155 = ~i6 & n154;
  assign n156 = i7 & n155;
  assign n157 = ~i2 & i3;
  assign n158 = ~i6 & n157;
  assign n159 = i7 & n158;
  assign n160 = ~i8 & n159;
  assign n161 = ~i9 & n160;
  assign n162 = ~i6 & n135;
  assign n163 = i7 & n162;
  assign n164 = ~i9 & n163;
  assign n165 = i2 & ~i3;
  assign n166 = i6 & n165;
  assign n167 = ~i8 & n166;
  assign n168 = ~i9 & n167;
  assign n169 = i6 & n154;
  assign n170 = ~i7 & n169;
  assign n171 = ~i9 & n82;
  assign n172 = i3 & n130;
  assign n173 = i6 & n172;
  assign n174 = i8 & n173;
  assign n175 = i6 & n157;
  assign n176 = ~i7 & n175;
  assign n177 = ~i8 & n176;
  assign n178 = ~i9 & n177;
  assign n179 = i2 & i3;
  assign n180 = ~i6 & n179;
  assign n181 = ~i7 & n180;
  assign n182 = ~i8 & n181;
  assign n183 = ~i9 & n182;
  assign n184 = ~i6 & n104;
  assign n185 = ~i7 & n184;
  assign n186 = ~i8 & n185;
  assign n187 = i3 & n146;
  assign n188 = ~i6 & n187;
  assign n189 = ~i7 & n188;
  assign n190 = ~i9 & n189;
  assign n191 = i6 & n179;
  assign n192 = i7 & n191;
  assign n193 = ~i8 & n192;
  assign n194 = ~i9 & n193;
  assign n195 = i6 & n187;
  assign n196 = i7 & n195;
  assign n197 = ~i9 & n196;
  assign n198 = ~i9 & n185;
  assign n199 = ~n38 & ~n42;
  assign n200 = ~n46 & n199;
  assign n201 = ~n50 & n200;
  assign n202 = ~n54 & n201;
  assign n203 = ~n59 & n202;
  assign n204 = ~n64 & n203;
  assign n205 = ~n68 & n204;
  assign n206 = ~n73 & n205;
  assign n207 = ~n74 & n206;
  assign n208 = ~n77 & n207;
  assign n209 = ~n80 & n208;
  assign n210 = ~n83 & n209;
  assign n211 = ~n84 & n210;
  assign n212 = ~n89 & n211;
  assign n213 = ~n94 & n212;
  assign n214 = ~n98 & n213;
  assign n215 = ~n100 & n214;
  assign n216 = ~n102 & n215;
  assign n217 = ~n107 & n216;
  assign n218 = ~n110 & n217;
  assign n219 = ~n111 & n218;
  assign n220 = ~n115 & n219;
  assign n221 = ~n119 & n220;
  assign n222 = ~n123 & n221;
  assign n223 = ~n126 & n222;
  assign n224 = ~n129 & n223;
  assign n225 = ~n134 & n224;
  assign n226 = ~n138 & n225;
  assign n227 = ~n141 & n226;
  assign n228 = ~n145 & n227;
  assign n229 = ~n149 & n228;
  assign n230 = ~n152 & n229;
  assign n231 = ~n153 & n230;
  assign n232 = ~n156 & n231;
  assign n233 = ~n161 & n232;
  assign n234 = ~n164 & n233;
  assign n235 = ~n168 & n234;
  assign n236 = ~n170 & n235;
  assign n237 = ~n171 & n236;
  assign n238 = ~n174 & n237;
  assign n239 = ~n178 & n238;
  assign n240 = ~n183 & n239;
  assign n241 = ~n186 & n240;
  assign n242 = ~n190 & n241;
  assign n243 = ~n194 & n242;
  assign n244 = ~n197 & n243;
  assign i10 = ~n198 & n244;
  assign n246 = i3 & n16;
  assign n247 = ~i7 & n246;
  assign n248 = i8 & n247;
  assign n249 = i0 & i3;
  assign n250 = ~i7 & n249;
  assign n251 = i9 & n250;
  assign n252 = i1 & i3;
  assign n253 = ~i7 & n252;
  assign n254 = i8 & n253;
  assign n255 = i9 & n254;
  assign n256 = i1 & ~i3;
  assign n257 = i7 & n256;
  assign n258 = i8 & n257;
  assign n259 = i9 & n258;
  assign n260 = n158 & ~i10;
  assign n261 = ~i0 & i3;
  assign n262 = i7 & n261;
  assign n263 = ~i9 & n262;
  assign n264 = ~i3 & n22;
  assign n265 = ~i7 & n264;
  assign n266 = n175 & i10;
  assign n267 = ~i0 & ~i3;
  assign n268 = ~i7 & n267;
  assign n269 = ~i9 & n268;
  assign n270 = n191 & ~i10;
  assign n271 = n180 & i10;
  assign n272 = ~i8 & n268;
  assign n273 = ~i1 & ~i3;
  assign n274 = ~i7 & n273;
  assign n275 = ~i9 & n274;
  assign n276 = ~i3 & ~i7;
  assign n277 = ~i8 & n276;
  assign n278 = ~i9 & n277;
  assign n279 = i0 & ~i3;
  assign n280 = i7 & n279;
  assign n281 = i9 & n280;
  assign n282 = ~i1 & i3;
  assign n283 = ~i7 & n282;
  assign n284 = ~i9 & n283;
  assign n285 = ~i3 & n16;
  assign n286 = i7 & n285;
  assign n287 = i8 & n286;
  assign n288 = i3 & n22;
  assign n289 = ~i7 & n288;
  assign n290 = ~i7 & n261;
  assign n291 = ~i9 & n290;
  assign n292 = i3 & ~i7;
  assign n293 = ~i8 & n292;
  assign n294 = ~i9 & n293;
  assign n295 = ~i8 & n290;
  assign n296 = ~n248 & ~n251;
  assign n297 = ~n255 & n296;
  assign n298 = ~n259 & n297;
  assign n299 = ~n260 & n298;
  assign n300 = ~n263 & n299;
  assign n301 = ~n265 & n300;
  assign n302 = ~n266 & n301;
  assign n303 = ~n269 & n302;
  assign n304 = ~n270 & n303;
  assign n305 = ~n270 & n304;
  assign n306 = ~n271 & n305;
  assign n307 = ~n272 & n306;
  assign n308 = ~n275 & n307;
  assign n309 = ~n278 & n308;
  assign n310 = ~n281 & n309;
  assign n311 = ~n284 & ~n310;
  assign n312 = ~n287 & ~n311;
  assign n313 = ~n260 & n312;
  assign n314 = ~n260 & n313;
  assign n315 = ~n260 & n314;
  assign n316 = ~n289 & ~n315;
  assign n317 = ~n291 & n316;
  assign n318 = ~n294 & n317;
  assign n319 = ~n295 & n318;
  assign n320 = ~n270 & ~n319;
  assign i11 = ~n270 & n320;
endmodule


