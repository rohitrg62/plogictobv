// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:27:17 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8, i9, i10, i11  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8, i9, i10, i11;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
    n27, n28, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
    n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
    n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
    n84, n85, n86, n87, n88, n89, n90, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
    n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
    n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466, n467;
  assign n13 = ~i0 & i1;
  assign n14 = i2 & n13;
  assign n15 = ~i3 & n14;
  assign n16 = i4 & n15;
  assign n17 = i5 & n16;
  assign n18 = i5 & ~i6;
  assign n19 = i5 & ~n18;
  assign n20 = i5 & i6;
  assign n21 = ~i7 & n20;
  assign n22 = ~i2 & n21;
  assign n23 = n19 & ~n22;
  assign n24 = i2 & n21;
  assign n25 = n23 & ~n24;
  assign n26 = i7 & n20;
  assign n27 = ~i4 & n26;
  assign n28 = n25 & ~n27;
  assign i11 = n17 | ~n28;
  assign n30 = i0 & ~i1;
  assign n31 = i2 & n30;
  assign n32 = ~i3 & n31;
  assign n33 = i4 & n32;
  assign n34 = ~i5 & n33;
  assign n35 = ~i5 & n16;
  assign n36 = i0 & i2;
  assign n37 = ~i3 & n36;
  assign n38 = ~i4 & n37;
  assign n39 = i5 & n38;
  assign n40 = ~i6 & n39;
  assign n41 = i7 & n40;
  assign n42 = i11 & n41;
  assign n43 = i5 & n15;
  assign n44 = i5 & n33;
  assign n45 = ~i6 & n44;
  assign n46 = ~i7 & n45;
  assign n47 = i11 & n46;
  assign n48 = i4 & n37;
  assign n49 = ~i5 & n48;
  assign n50 = ~i7 & n49;
  assign n51 = ~i4 & n32;
  assign n52 = i5 & n51;
  assign n53 = ~i0 & ~i1;
  assign n54 = i2 & n53;
  assign n55 = i3 & n54;
  assign n56 = i4 & n55;
  assign n57 = ~i5 & n56;
  assign n58 = ~i7 & n57;
  assign n59 = i7 & n39;
  assign n60 = i11 & n59;
  assign n61 = ~i4 & n36;
  assign n62 = i5 & n61;
  assign n63 = i6 & n62;
  assign n64 = i7 & n63;
  assign n65 = i11 & n64;
  assign n66 = ~i4 & n55;
  assign n67 = i5 & n66;
  assign n68 = i6 & n67;
  assign n69 = i7 & n68;
  assign n70 = i11 & n69;
  assign n71 = ~i4 & n14;
  assign n72 = i5 & n71;
  assign n73 = i6 & n72;
  assign n74 = i7 & n73;
  assign n75 = i11 & n74;
  assign n76 = ~i6 & i11;
  assign n77 = i11 & ~n76;
  assign n78 = i6 & i11;
  assign n79 = n77 & ~n78;
  assign n80 = ~n34 & ~n79;
  assign n81 = ~n35 & n80;
  assign n82 = ~n42 & n81;
  assign n83 = ~n43 & n82;
  assign n84 = ~n47 & n83;
  assign n85 = ~n50 & n84;
  assign n86 = ~n52 & n85;
  assign n87 = ~n58 & n86;
  assign n88 = ~n60 & n87;
  assign n89 = ~n65 & n88;
  assign n90 = ~n70 & n89;
  assign i8 = ~n75 & n90;
  assign n92 = n41 & ~i8;
  assign n93 = i11 & n92;
  assign n94 = i4 & n14;
  assign n95 = i5 & n94;
  assign n96 = i7 & n95;
  assign n97 = i8 & n96;
  assign n98 = i1 & i2;
  assign n99 = ~i3 & n98;
  assign n100 = ~i4 & n99;
  assign n101 = i5 & n100;
  assign n102 = ~i6 & n101;
  assign n103 = i7 & n102;
  assign n104 = ~i8 & n103;
  assign n105 = i11 & n104;
  assign n106 = n17 & ~i8;
  assign n107 = i4 & n36;
  assign n108 = i5 & n107;
  assign n109 = ~i6 & n108;
  assign n110 = ~i7 & n109;
  assign n111 = ~i8 & n110;
  assign n112 = i11 & n111;
  assign n113 = ~i4 & n15;
  assign n114 = i5 & n113;
  assign n115 = ~i2 & n13;
  assign n116 = ~i3 & n115;
  assign n117 = ~i4 & n116;
  assign n118 = i5 & n117;
  assign n119 = i6 & n118;
  assign n120 = i7 & n119;
  assign n121 = i8 & n120;
  assign n122 = i11 & n121;
  assign n123 = ~i2 & n53;
  assign n124 = ~i3 & n123;
  assign n125 = ~i4 & n124;
  assign n126 = i5 & n125;
  assign n127 = i6 & n126;
  assign n128 = i7 & n127;
  assign n129 = i8 & n128;
  assign n130 = i11 & n129;
  assign n131 = i4 & n124;
  assign n132 = ~i5 & n131;
  assign n133 = i6 & n132;
  assign n134 = i7 & n133;
  assign n135 = i8 & n134;
  assign n136 = i4 & n116;
  assign n137 = ~i5 & n136;
  assign n138 = i6 & n137;
  assign n139 = i7 & n138;
  assign n140 = i8 & n139;
  assign n141 = ~i7 & n39;
  assign n142 = i5 & n56;
  assign n143 = i7 & n142;
  assign n144 = i8 & n143;
  assign n145 = ~i7 & n44;
  assign n146 = i8 & n145;
  assign n147 = ~i2 & n30;
  assign n148 = ~i3 & n147;
  assign n149 = i4 & n148;
  assign n150 = ~i5 & n149;
  assign n151 = i6 & n150;
  assign n152 = i7 & n151;
  assign n153 = i8 & n152;
  assign n154 = i4 & n98;
  assign n155 = ~i5 & n154;
  assign n156 = i6 & n155;
  assign n157 = i7 & n156;
  assign n158 = i8 & n157;
  assign n159 = ~i7 & n72;
  assign n160 = i8 & n159;
  assign n161 = ~i7 & n67;
  assign n162 = i0 & ~i2;
  assign n163 = ~i3 & n162;
  assign n164 = ~i4 & n163;
  assign n165 = i5 & n164;
  assign n166 = i6 & n165;
  assign n167 = i7 & n166;
  assign n168 = i8 & n167;
  assign n169 = i11 & n168;
  assign n170 = ~i4 & n31;
  assign n171 = i5 & n170;
  assign n172 = ~i7 & n171;
  assign n173 = i8 & n172;
  assign n174 = ~i5 & n107;
  assign n175 = i6 & n174;
  assign n176 = i7 & n175;
  assign n177 = i8 & n176;
  assign n178 = i6 & n57;
  assign n179 = i7 & n178;
  assign n180 = i8 & n179;
  assign n181 = ~i4 & ~i5;
  assign n182 = i4 & ~i5;
  assign n183 = ~i6 & n182;
  assign n184 = ~n181 & ~n183;
  assign n185 = i6 & n182;
  assign n186 = n184 & ~n185;
  assign n187 = i5 & ~i7;
  assign n188 = n186 & ~n187;
  assign n189 = i5 & i7;
  assign n190 = ~i11 & n189;
  assign n191 = i0 & n190;
  assign n192 = n188 & ~n191;
  assign n193 = i11 & n189;
  assign n194 = n192 & ~n193;
  assign n195 = ~n93 & ~n194;
  assign n196 = ~n97 & ~n195;
  assign n197 = ~n105 & ~n196;
  assign n198 = ~n106 & n197;
  assign n199 = ~n112 & n198;
  assign n200 = ~n114 & n199;
  assign n201 = ~n122 & n200;
  assign n202 = ~n130 & n201;
  assign n203 = ~n135 & n202;
  assign n204 = ~n140 & n203;
  assign n205 = ~n141 & n204;
  assign n206 = ~n144 & ~n205;
  assign n207 = ~n146 & ~n206;
  assign n208 = ~n153 & n207;
  assign n209 = ~n158 & n208;
  assign n210 = ~n160 & n209;
  assign n211 = ~n161 & n210;
  assign n212 = ~n169 & n211;
  assign n213 = ~n173 & n212;
  assign n214 = ~n177 & n213;
  assign i10 = ~n180 & n214;
  assign n216 = ~i4 & n123;
  assign n217 = ~i5 & n216;
  assign n218 = i6 & n217;
  assign n219 = i7 & n218;
  assign n220 = i8 & n219;
  assign n221 = i4 & n31;
  assign n222 = ~i5 & n221;
  assign n223 = i7 & n222;
  assign n224 = ~i8 & n223;
  assign n225 = ~i5 & n94;
  assign n226 = i7 & n225;
  assign n227 = ~i8 & n226;
  assign n228 = n59 & ~i10;
  assign n229 = ~i5 & n66;
  assign n230 = i7 & n229;
  assign n231 = ~i5 & n38;
  assign n232 = i7 & n231;
  assign n233 = ~i5 & n100;
  assign n234 = i7 & n233;
  assign n235 = ~i7 & n142;
  assign n236 = i8 & n235;
  assign n237 = i10 & n236;
  assign n238 = i7 & n72;
  assign n239 = ~i10 & n238;
  assign n240 = i5 & n154;
  assign n241 = i7 & n240;
  assign n242 = ~i8 & n241;
  assign n243 = ~i10 & n242;
  assign n244 = n33 & ~i8;
  assign n245 = ~i5 & n164;
  assign n246 = i6 & n245;
  assign n247 = i7 & n246;
  assign n248 = i8 & n247;
  assign n249 = i1 & ~i2;
  assign n250 = ~i3 & n249;
  assign n251 = ~i4 & n250;
  assign n252 = ~i5 & n251;
  assign n253 = i6 & n252;
  assign n254 = i7 & n253;
  assign n255 = i8 & n254;
  assign n256 = ~i4 & n98;
  assign n257 = i5 & n256;
  assign n258 = i6 & n257;
  assign n259 = ~i8 & n258;
  assign n260 = ~i10 & n259;
  assign n261 = i11 & n260;
  assign n262 = ~i7 & n175;
  assign n263 = ~i8 & n262;
  assign n264 = i10 & n263;
  assign n265 = ~i7 & n133;
  assign n266 = i10 & n265;
  assign n267 = ~i7 & n151;
  assign n268 = i10 & n267;
  assign n269 = ~i7 & n138;
  assign n270 = i10 & n269;
  assign n271 = ~i7 & n62;
  assign n272 = i8 & n271;
  assign n273 = i10 & n272;
  assign n274 = n39 & i8;
  assign n275 = i4 & n163;
  assign n276 = ~i5 & n275;
  assign n277 = i6 & n276;
  assign n278 = ~i7 & n277;
  assign n279 = i8 & n278;
  assign n280 = i10 & n279;
  assign n281 = i5 & n48;
  assign n282 = ~i7 & n281;
  assign n283 = i8 & n282;
  assign n284 = i10 & n283;
  assign n285 = n44 & i8;
  assign n286 = ~i5 & n61;
  assign n287 = i6 & n286;
  assign n288 = i7 & n287;
  assign n289 = i8 & n288;
  assign n290 = i2 & i3;
  assign n291 = i4 & n290;
  assign n292 = ~i5 & n291;
  assign n293 = i6 & n292;
  assign n294 = ~i7 & n293;
  assign n295 = ~i8 & n294;
  assign n296 = i10 & n295;
  assign n297 = i3 & n123;
  assign n298 = ~i4 & n297;
  assign n299 = i5 & n298;
  assign n300 = i6 & n299;
  assign n301 = ~i7 & n300;
  assign n302 = i10 & n301;
  assign n303 = i11 & n302;
  assign n304 = ~i7 & n63;
  assign n305 = ~i10 & n304;
  assign n306 = i11 & n305;
  assign n307 = i6 & n108;
  assign n308 = ~i7 & n307;
  assign n309 = i8 & n308;
  assign n310 = i10 & n309;
  assign n311 = i11 & n310;
  assign n312 = n39 & i10;
  assign n313 = i4 & n297;
  assign n314 = ~i5 & n313;
  assign n315 = i6 & n314;
  assign n316 = ~i7 & n315;
  assign n317 = i8 & n316;
  assign n318 = i10 & n317;
  assign n319 = ~i7 & n127;
  assign n320 = i11 & n319;
  assign n321 = ~i5 & n256;
  assign n322 = i6 & n321;
  assign n323 = i7 & n322;
  assign n324 = i8 & n323;
  assign n325 = i4 & n115;
  assign n326 = ~i5 & n325;
  assign n327 = i6 & n326;
  assign n328 = ~i7 & n327;
  assign n329 = i8 & n328;
  assign n330 = i10 & n329;
  assign n331 = i5 & n251;
  assign n332 = i6 & n331;
  assign n333 = ~i7 & n332;
  assign n334 = i8 & n333;
  assign n335 = i11 & n334;
  assign n336 = i4 & n147;
  assign n337 = ~i5 & n336;
  assign n338 = i6 & n337;
  assign n339 = ~i7 & n338;
  assign n340 = i8 & n339;
  assign n341 = i10 & n340;
  assign n342 = ~i7 & n225;
  assign n343 = i8 & n342;
  assign n344 = ~i7 & n222;
  assign n345 = i8 & n344;
  assign n346 = ~i4 & n249;
  assign n347 = i5 & n346;
  assign n348 = i6 & n347;
  assign n349 = ~i7 & n348;
  assign n350 = i8 & n349;
  assign n351 = i10 & n350;
  assign n352 = i11 & n351;
  assign n353 = ~i4 & n148;
  assign n354 = i5 & n353;
  assign n355 = i6 & n354;
  assign n356 = ~i7 & n355;
  assign n357 = i8 & n356;
  assign n358 = i11 & n357;
  assign n359 = i5 & n131;
  assign n360 = i6 & n359;
  assign n361 = ~i7 & n360;
  assign n362 = i8 & n361;
  assign n363 = i10 & n362;
  assign n364 = i11 & n363;
  assign n365 = ~i4 & n147;
  assign n366 = i5 & n365;
  assign n367 = i6 & n366;
  assign n368 = ~i7 & n367;
  assign n369 = i8 & n368;
  assign n370 = i10 & n369;
  assign n371 = i11 & n370;
  assign n372 = ~i7 & n95;
  assign n373 = i8 & n372;
  assign n374 = i10 & n373;
  assign n375 = i5 & n325;
  assign n376 = i6 & n375;
  assign n377 = ~i7 & n376;
  assign n378 = i8 & n377;
  assign n379 = i10 & n378;
  assign n380 = i11 & n379;
  assign n381 = i5 & n275;
  assign n382 = i6 & n381;
  assign n383 = ~i7 & n382;
  assign n384 = i8 & n383;
  assign n385 = i10 & n384;
  assign n386 = i11 & n385;
  assign n387 = i5 & n313;
  assign n388 = i6 & n387;
  assign n389 = ~i7 & n388;
  assign n390 = i8 & n389;
  assign n391 = i10 & n390;
  assign n392 = i11 & n391;
  assign n393 = ~i7 & n258;
  assign n394 = ~i10 & n393;
  assign n395 = i11 & n394;
  assign n396 = ~i4 & n290;
  assign n397 = i5 & n396;
  assign n398 = i6 & n397;
  assign n399 = ~i7 & n398;
  assign n400 = ~i10 & n399;
  assign n401 = i11 & n400;
  assign n402 = i10 & n262;
  assign n403 = ~i4 & ~i10;
  assign n404 = ~i2 & n403;
  assign n405 = i2 & n403;
  assign n406 = ~i7 & n405;
  assign n407 = ~n404 & ~n406;
  assign n408 = i4 & ~i10;
  assign n409 = ~i8 & n408;
  assign n410 = ~i1 & n409;
  assign n411 = n407 & ~n410;
  assign n412 = i8 & n408;
  assign n413 = n411 & ~n412;
  assign n414 = ~i6 & i10;
  assign n415 = n413 & ~n414;
  assign n416 = i6 & i10;
  assign n417 = n415 & ~n416;
  assign n418 = ~n220 & ~n417;
  assign n419 = ~n224 & n418;
  assign n420 = ~n227 & n419;
  assign n421 = ~n228 & n420;
  assign n422 = ~n230 & n421;
  assign n423 = ~n232 & n422;
  assign n424 = ~n234 & n423;
  assign n425 = ~n237 & n424;
  assign n426 = ~n34 & n425;
  assign n427 = ~n239 & n426;
  assign n428 = ~n243 & n427;
  assign n429 = ~n244 & n428;
  assign n430 = ~n248 & n429;
  assign n431 = ~n255 & n430;
  assign n432 = ~n16 & n431;
  assign n433 = ~n261 & n432;
  assign n434 = ~n43 & n433;
  assign n435 = ~n264 & n434;
  assign n436 = ~n266 & n435;
  assign n437 = ~n268 & n436;
  assign n438 = ~n270 & n437;
  assign n439 = ~n273 & n438;
  assign n440 = ~n274 & n439;
  assign n441 = ~n280 & n440;
  assign n442 = ~n284 & n441;
  assign n443 = ~n285 & ~n442;
  assign n444 = ~n289 & ~n443;
  assign n445 = ~n296 & n444;
  assign n446 = ~n303 & n445;
  assign n447 = ~n306 & n446;
  assign n448 = ~n311 & n447;
  assign n449 = ~n312 & ~n448;
  assign n450 = ~n318 & ~n449;
  assign n451 = ~n320 & n450;
  assign n452 = ~n324 & n451;
  assign n453 = ~n330 & n452;
  assign n454 = ~n335 & n453;
  assign n455 = ~n341 & n454;
  assign n456 = ~n343 & n455;
  assign n457 = ~n345 & n456;
  assign n458 = ~n352 & n457;
  assign n459 = ~n358 & n458;
  assign n460 = ~n364 & n459;
  assign n461 = ~n371 & n460;
  assign n462 = ~n374 & n461;
  assign n463 = ~n380 & n462;
  assign n464 = ~n386 & n463;
  assign n465 = ~n392 & n464;
  assign n466 = ~n395 & n465;
  assign n467 = ~n401 & n466;
  assign i9 = ~n402 & n467;
endmodule


