// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:27:42 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8, i9, i10, i11  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8, i9, i10, i11;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n25, n26, n27,
    n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
    n42, n43, n44, n45, n46, n47, n48, n49, n50, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
    n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n111,
    n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
    n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253;
  assign n13 = ~i1 & ~i5;
  assign n14 = ~i7 & n13;
  assign n15 = ~i6 & n14;
  assign n16 = i4 & n15;
  assign n17 = ~i3 & n16;
  assign n18 = i6 & n14;
  assign n19 = ~n17 & ~n18;
  assign n20 = i7 & n13;
  assign n21 = n19 & ~n20;
  assign n22 = ~i1 & i5;
  assign n23 = n21 & ~n22;
  assign i8 = i1 | ~n23;
  assign n25 = i2 & i3;
  assign n26 = ~i4 & n25;
  assign n27 = ~i5 & n26;
  assign n28 = ~i6 & n27;
  assign n29 = ~i7 & n28;
  assign n30 = i8 & n29;
  assign n31 = ~i0 & ~i1;
  assign n32 = ~i2 & n31;
  assign n33 = ~i3 & n32;
  assign n34 = ~i6 & n33;
  assign n35 = ~i7 & n34;
  assign n36 = ~i4 & n33;
  assign n37 = ~i5 & n36;
  assign n38 = ~i6 & n37;
  assign n39 = i8 & n38;
  assign n40 = i2 & n31;
  assign n41 = ~i3 & n40;
  assign n42 = ~i4 & n41;
  assign n43 = ~i5 & n42;
  assign n44 = ~i6 & n43;
  assign n45 = i8 & n44;
  assign n46 = ~i2 & ~i7;
  assign n47 = ~i7 & ~n46;
  assign n48 = ~n30 & n47;
  assign n49 = ~n35 & ~n48;
  assign n50 = ~n39 & n49;
  assign i10 = ~n45 & n50;
  assign n52 = i2 & ~i4;
  assign n53 = ~i5 & n52;
  assign n54 = ~i6 & n53;
  assign n55 = ~i7 & n54;
  assign n56 = i8 & n55;
  assign n57 = i8 & n37;
  assign n58 = i10 & n57;
  assign n59 = i0 & ~i2;
  assign n60 = i3 & n59;
  assign n61 = ~i4 & n60;
  assign n62 = ~i5 & n61;
  assign n63 = ~i6 & n62;
  assign n64 = ~i7 & n63;
  assign n65 = i8 & n64;
  assign n66 = i10 & n65;
  assign n67 = ~i7 & n33;
  assign n68 = i10 & n67;
  assign n69 = i0 & ~i1;
  assign n70 = i2 & n69;
  assign n71 = i3 & n70;
  assign n72 = ~i4 & n71;
  assign n73 = ~i5 & n72;
  assign n74 = ~i7 & n73;
  assign n75 = i8 & n74;
  assign n76 = ~i10 & n75;
  assign n77 = i3 & n40;
  assign n78 = ~i4 & n77;
  assign n79 = ~i5 & n78;
  assign n80 = ~i7 & n79;
  assign n81 = i8 & n80;
  assign n82 = ~i10 & n81;
  assign n83 = ~i7 & n27;
  assign n84 = i8 & n83;
  assign n85 = ~i10 & n84;
  assign n86 = i6 & ~i10;
  assign n87 = ~i6 & ~i10;
  assign n88 = ~i3 & n87;
  assign n89 = ~i1 & n88;
  assign n90 = i2 & n89;
  assign n91 = ~i0 & n90;
  assign n92 = i1 & n88;
  assign n93 = ~n91 & ~n92;
  assign n94 = i3 & n87;
  assign n95 = ~i2 & n94;
  assign n96 = i8 & n95;
  assign n97 = n93 & ~n96;
  assign n98 = ~n86 & n97;
  assign n99 = ~i4 & i10;
  assign n100 = n98 & ~n99;
  assign n101 = i4 & i10;
  assign n102 = n100 & ~n101;
  assign n103 = ~n56 & n102;
  assign n104 = ~n34 & ~n103;
  assign n105 = ~n58 & n104;
  assign n106 = ~n66 & n105;
  assign n107 = ~n68 & n106;
  assign n108 = ~n76 & n107;
  assign n109 = ~n82 & n108;
  assign i9 = ~n85 & n109;
  assign n111 = ~i0 & i2;
  assign n112 = ~i5 & n111;
  assign n113 = ~i6 & n112;
  assign n114 = ~i7 & n113;
  assign n115 = i8 & n114;
  assign n116 = ~i9 & n115;
  assign n117 = ~i5 & n70;
  assign n118 = ~i6 & n117;
  assign n119 = ~i7 & n118;
  assign n120 = i8 & n119;
  assign n121 = ~i9 & n120;
  assign n122 = i0 & i2;
  assign n123 = ~i5 & n122;
  assign n124 = ~i6 & n123;
  assign n125 = ~i7 & n124;
  assign n126 = i8 & n125;
  assign n127 = ~i9 & n126;
  assign n128 = ~i6 & n36;
  assign n129 = i10 & n128;
  assign n130 = ~i5 & n33;
  assign n131 = ~i6 & n130;
  assign n132 = i8 & n131;
  assign n133 = i10 & n132;
  assign n134 = ~i3 & n70;
  assign n135 = ~i4 & n134;
  assign n136 = ~i5 & n135;
  assign n137 = ~i6 & n136;
  assign n138 = i8 & n137;
  assign n139 = i9 & n138;
  assign n140 = i10 & n139;
  assign n141 = ~i4 & n111;
  assign n142 = ~i6 & n141;
  assign n143 = ~i7 & n142;
  assign n144 = i8 & n143;
  assign n145 = ~i4 & n31;
  assign n146 = ~i6 & n145;
  assign n147 = ~i7 & n146;
  assign n148 = ~i6 & n42;
  assign n149 = i9 & n148;
  assign n150 = i10 & n149;
  assign n151 = ~i5 & n41;
  assign n152 = ~i6 & n151;
  assign n153 = i8 & n152;
  assign n154 = i9 & n153;
  assign n155 = i10 & n154;
  assign n156 = i8 & n130;
  assign n157 = i9 & n156;
  assign n158 = i10 & n157;
  assign n159 = n36 & i9;
  assign n160 = i10 & n159;
  assign n161 = ~i7 & n131;
  assign n162 = i8 & n161;
  assign n163 = ~i5 & n31;
  assign n164 = ~i6 & n163;
  assign n165 = ~i7 & n164;
  assign n166 = i8 & n165;
  assign n167 = ~i5 & n77;
  assign n168 = ~i7 & n167;
  assign n169 = i8 & n168;
  assign n170 = i9 & n169;
  assign n171 = ~i10 & n170;
  assign n172 = ~i2 & n69;
  assign n173 = i3 & n172;
  assign n174 = ~i4 & n173;
  assign n175 = ~i6 & n174;
  assign n176 = ~i7 & n175;
  assign n177 = i9 & n176;
  assign n178 = i10 & n177;
  assign n179 = ~i0 & i1;
  assign n180 = i2 & n179;
  assign n181 = ~i3 & n180;
  assign n182 = ~i4 & n181;
  assign n183 = ~i6 & n182;
  assign n184 = i8 & n183;
  assign n185 = i10 & n184;
  assign n186 = i0 & i1;
  assign n187 = i2 & n186;
  assign n188 = ~i6 & n187;
  assign n189 = i9 & n188;
  assign n190 = ~i10 & n189;
  assign n191 = i3 & n111;
  assign n192 = ~i5 & n191;
  assign n193 = ~i7 & n192;
  assign n194 = i8 & n193;
  assign n195 = i9 & n194;
  assign n196 = ~i10 & n195;
  assign n197 = ~i7 & n78;
  assign n198 = i9 & n197;
  assign n199 = ~i10 & n198;
  assign n200 = ~i7 & n72;
  assign n201 = i9 & n200;
  assign n202 = ~i10 & n201;
  assign n203 = ~i5 & n71;
  assign n204 = ~i7 & n203;
  assign n205 = i8 & n204;
  assign n206 = i9 & n205;
  assign n207 = ~i10 & n206;
  assign n208 = i3 & n187;
  assign n209 = ~i4 & n208;
  assign n210 = ~i7 & n209;
  assign n211 = i8 & n210;
  assign n212 = i9 & n211;
  assign n213 = ~i10 & n212;
  assign n214 = ~i4 & n191;
  assign n215 = ~i7 & n214;
  assign n216 = i8 & n215;
  assign n217 = i9 & n216;
  assign n218 = ~i10 & n217;
  assign n219 = ~i5 & n208;
  assign n220 = ~i7 & n219;
  assign n221 = i8 & n220;
  assign n222 = i9 & n221;
  assign n223 = ~i10 & n222;
  assign n224 = ~i4 & ~i6;
  assign n225 = i8 & n224;
  assign n226 = i10 & n225;
  assign n227 = i4 & ~i6;
  assign n228 = ~n226 & ~n227;
  assign n229 = ~i6 & n228;
  assign n230 = ~n116 & ~n229;
  assign n231 = ~n121 & n230;
  assign n232 = ~n127 & n231;
  assign n233 = ~n129 & n232;
  assign n234 = ~n133 & n233;
  assign n235 = ~n140 & n234;
  assign n236 = ~n144 & n235;
  assign n237 = ~n147 & n236;
  assign n238 = ~n150 & n237;
  assign n239 = ~n155 & n238;
  assign n240 = ~n158 & n239;
  assign n241 = ~n160 & n240;
  assign n242 = ~n162 & n241;
  assign n243 = ~n166 & n242;
  assign n244 = ~n171 & n243;
  assign n245 = ~n178 & n244;
  assign n246 = ~n185 & n245;
  assign n247 = ~n190 & ~n246;
  assign n248 = ~n196 & ~n247;
  assign n249 = ~n199 & n248;
  assign n250 = ~n202 & n249;
  assign n251 = ~n207 & n250;
  assign n252 = ~n213 & n251;
  assign n253 = ~n218 & n252;
  assign i11 = ~n223 & n253;
endmodule


