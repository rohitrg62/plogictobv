// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:26:50 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8, i9, i10, i11  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8, i9, i10, i11;
  assign i8 = 1'b0;
  assign i9 = 1'b0;
  assign i10 = 1'b1;
  assign i11 = 1'b0;
endmodule


