// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:26:55 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8, i9, i10, i11  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8, i9, i10, i11;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
    n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
    n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n55,
    n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
    n84, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n152, n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320;
  assign n13 = ~i0 & ~i1;
  assign n14 = ~i3 & n13;
  assign n15 = ~i4 & n14;
  assign n16 = ~i5 & n15;
  assign n17 = ~i6 & n16;
  assign n18 = ~i7 & n17;
  assign n19 = i0 & ~i1;
  assign n20 = i2 & n19;
  assign n21 = ~i3 & n20;
  assign n22 = i4 & n21;
  assign n23 = i5 & n22;
  assign n24 = i6 & n23;
  assign n25 = ~i4 & n13;
  assign n26 = ~i5 & n25;
  assign n27 = ~i6 & n26;
  assign n28 = ~i7 & n27;
  assign n29 = ~i0 & ~i4;
  assign n30 = ~i5 & n29;
  assign n31 = ~i6 & n30;
  assign n32 = ~i7 & n31;
  assign n33 = ~i0 & ~i6;
  assign n34 = i2 & n33;
  assign n35 = ~i3 & n34;
  assign n36 = i3 & n34;
  assign n37 = ~n35 & ~n36;
  assign n38 = i0 & ~i5;
  assign n39 = n37 & ~n38;
  assign n40 = i0 & i5;
  assign n41 = ~i6 & n40;
  assign n42 = i4 & n41;
  assign n43 = ~i3 & n42;
  assign n44 = n39 & ~n43;
  assign n45 = i6 & n40;
  assign n46 = ~i7 & n45;
  assign n47 = ~i2 & n46;
  assign n48 = n44 & ~n47;
  assign n49 = i7 & n45;
  assign n50 = n48 & ~n49;
  assign n51 = ~n18 & ~n50;
  assign n52 = ~n24 & ~n51;
  assign n53 = ~n28 & ~n52;
  assign i9 = ~n32 & n53;
  assign n55 = ~i2 & n13;
  assign n56 = i4 & n55;
  assign n57 = i5 & n56;
  assign n58 = i7 & n57;
  assign n59 = ~i9 & n58;
  assign n60 = ~i5 & n56;
  assign n61 = i7 & n60;
  assign n62 = ~i1 & ~i2;
  assign n63 = ~i4 & n62;
  assign n64 = ~i5 & n63;
  assign n65 = ~i6 & n64;
  assign n66 = ~i7 & n65;
  assign n67 = ~i1 & ~i4;
  assign n68 = ~i5 & n67;
  assign n69 = ~i6 & n68;
  assign n70 = ~i7 & n69;
  assign n71 = i1 & ~i5;
  assign n72 = ~i1 & ~i6;
  assign n73 = ~i2 & n72;
  assign n74 = i3 & n73;
  assign n75 = i2 & n72;
  assign n76 = ~n74 & ~n75;
  assign n77 = ~n71 & n76;
  assign n78 = i1 & i5;
  assign n79 = n77 & ~n78;
  assign n80 = ~n18 & ~n79;
  assign n81 = ~n59 & n80;
  assign n82 = ~n61 & n81;
  assign n83 = ~n28 & n82;
  assign n84 = ~n66 & n83;
  assign i11 = ~n70 & n84;
  assign n86 = ~i2 & n19;
  assign n87 = ~i3 & n86;
  assign n88 = i5 & n87;
  assign n89 = i7 & n88;
  assign n90 = ~i9 & n89;
  assign n91 = ~i11 & n90;
  assign n92 = i0 & ~i2;
  assign n93 = ~i3 & n92;
  assign n94 = ~i4 & n93;
  assign n95 = i5 & n94;
  assign n96 = i7 & n95;
  assign n97 = ~i9 & n96;
  assign n98 = i11 & n97;
  assign n99 = i2 & n13;
  assign n100 = ~i3 & n99;
  assign n101 = i5 & n100;
  assign n102 = i6 & n101;
  assign n103 = ~i7 & n102;
  assign n104 = ~i1 & i2;
  assign n105 = ~i3 & n104;
  assign n106 = i4 & n105;
  assign n107 = i5 & n106;
  assign n108 = i6 & n107;
  assign n109 = ~i7 & n108;
  assign n110 = i4 & n87;
  assign n111 = i5 & n110;
  assign n112 = i7 & n111;
  assign n113 = i9 & n112;
  assign n114 = ~i11 & n113;
  assign n115 = i3 & n55;
  assign n116 = ~i4 & n115;
  assign n117 = i5 & n116;
  assign n118 = i7 & n117;
  assign n119 = ~i9 & n118;
  assign n120 = i11 & n119;
  assign n121 = i0 & i1;
  assign n122 = ~i2 & n121;
  assign n123 = ~i3 & n122;
  assign n124 = i4 & n123;
  assign n125 = i5 & n124;
  assign n126 = i7 & n125;
  assign n127 = i9 & n126;
  assign n128 = i11 & n127;
  assign n129 = ~i3 & ~i6;
  assign n130 = i4 & n129;
  assign n131 = i9 & n130;
  assign n132 = ~i3 & i6;
  assign n133 = i2 & n132;
  assign n134 = ~i7 & n133;
  assign n135 = ~i9 & n134;
  assign n136 = ~i0 & n135;
  assign n137 = ~i4 & n136;
  assign n138 = ~n131 & ~n137;
  assign n139 = i0 & n135;
  assign n140 = n138 & ~n139;
  assign n141 = i3 & ~i11;
  assign n142 = n140 & ~n141;
  assign n143 = i3 & i11;
  assign n144 = n142 & ~n143;
  assign n145 = ~n91 & n144;
  assign n146 = ~n98 & n145;
  assign n147 = ~n103 & ~n146;
  assign n148 = ~n109 & n147;
  assign n149 = ~n114 & n148;
  assign n150 = ~n120 & n149;
  assign i10 = ~n128 & n150;
  assign n152 = ~i4 & n100;
  assign n153 = ~i5 & n152;
  assign n154 = ~i6 & n153;
  assign n155 = ~i7 & n154;
  assign n156 = ~i2 & i4;
  assign n157 = ~i5 & n156;
  assign n158 = i6 & n157;
  assign n159 = ~i9 & n158;
  assign n160 = ~i10 & n159;
  assign n161 = i1 & ~i2;
  assign n162 = ~i4 & n161;
  assign n163 = i5 & n162;
  assign n164 = i6 & n163;
  assign n165 = ~i7 & n164;
  assign n166 = i11 & n165;
  assign n167 = ~i2 & i5;
  assign n168 = i6 & n167;
  assign n169 = ~i9 & n168;
  assign n170 = ~i10 & n169;
  assign n171 = ~i11 & n170;
  assign n172 = ~i2 & ~i3;
  assign n173 = ~i4 & n172;
  assign n174 = i5 & n173;
  assign n175 = ~i6 & n174;
  assign n176 = i7 & n175;
  assign n177 = ~i9 & n176;
  assign n178 = ~i10 & n177;
  assign n179 = i11 & n178;
  assign n180 = ~i6 & n57;
  assign n181 = i7 & n180;
  assign n182 = ~i9 & n181;
  assign n183 = ~i11 & n182;
  assign n184 = ~i0 & ~i2;
  assign n185 = i3 & n184;
  assign n186 = i4 & n185;
  assign n187 = ~i5 & n186;
  assign n188 = ~i6 & n187;
  assign n189 = i7 & n188;
  assign n190 = ~i9 & n189;
  assign n191 = i10 & n190;
  assign n192 = ~i4 & n92;
  assign n193 = i5 & n192;
  assign n194 = i6 & n193;
  assign n195 = ~i7 & n194;
  assign n196 = i9 & n195;
  assign n197 = ~i11 & n196;
  assign n198 = i4 & n184;
  assign n199 = i5 & n198;
  assign n200 = ~i6 & n199;
  assign n201 = i7 & n200;
  assign n202 = ~i9 & n201;
  assign n203 = i11 & n202;
  assign n204 = ~i4 & n99;
  assign n205 = ~i5 & n204;
  assign n206 = ~i6 & n205;
  assign n207 = ~i7 & n206;
  assign n208 = i6 & n156;
  assign n209 = ~i9 & n208;
  assign n210 = ~i10 & n209;
  assign n211 = ~i0 & i1;
  assign n212 = ~i2 & n211;
  assign n213 = ~i3 & n212;
  assign n214 = i4 & n213;
  assign n215 = i5 & n214;
  assign n216 = ~i6 & n215;
  assign n217 = ~i7 & n216;
  assign n218 = ~i9 & n217;
  assign n219 = ~i10 & n218;
  assign n220 = i11 & n219;
  assign n221 = ~i3 & n184;
  assign n222 = i4 & n221;
  assign n223 = i5 & n222;
  assign n224 = ~i6 & n223;
  assign n225 = ~i7 & n224;
  assign n226 = ~i9 & n225;
  assign n227 = ~i10 & n226;
  assign n228 = ~i11 & n227;
  assign n229 = ~i3 & n62;
  assign n230 = i4 & n229;
  assign n231 = i5 & n230;
  assign n232 = ~i6 & n231;
  assign n233 = i7 & n232;
  assign n234 = ~i10 & n233;
  assign n235 = ~i11 & n234;
  assign n236 = ~i5 & n222;
  assign n237 = ~i6 & n236;
  assign n238 = i7 & n237;
  assign n239 = ~i9 & n238;
  assign n240 = ~i10 & n239;
  assign n241 = i4 & n92;
  assign n242 = ~i5 & n241;
  assign n243 = i6 & n242;
  assign n244 = ~i7 & n243;
  assign n245 = i9 & n244;
  assign n246 = i5 & n156;
  assign n247 = i6 & n246;
  assign n248 = ~i10 & n247;
  assign n249 = ~i11 & n248;
  assign n250 = i2 & ~i4;
  assign n251 = ~i5 & n250;
  assign n252 = ~i6 & n251;
  assign n253 = ~i7 & n252;
  assign n254 = ~i3 & n55;
  assign n255 = ~i4 & n254;
  assign n256 = i5 & n255;
  assign n257 = ~i6 & n256;
  assign n258 = i7 & n257;
  assign n259 = ~i9 & n258;
  assign n260 = ~i10 & n259;
  assign n261 = ~i11 & n260;
  assign n262 = i6 & n241;
  assign n263 = ~i7 & n262;
  assign n264 = i9 & n263;
  assign n265 = i11 & n264;
  assign n266 = ~i3 & n161;
  assign n267 = i4 & n266;
  assign n268 = i5 & n267;
  assign n269 = ~i6 & n268;
  assign n270 = i7 & n269;
  assign n271 = ~i10 & n270;
  assign n272 = i11 & n271;
  assign n273 = ~i2 & ~i6;
  assign n274 = ~i5 & n273;
  assign n275 = ~i7 & n274;
  assign n276 = i4 & n275;
  assign n277 = ~i3 & n276;
  assign n278 = ~i9 & n277;
  assign n279 = i3 & n276;
  assign n280 = ~n278 & ~n279;
  assign n281 = i7 & n274;
  assign n282 = n280 & ~n281;
  assign n283 = i5 & n273;
  assign n284 = n282 & ~n283;
  assign n285 = ~i2 & i6;
  assign n286 = ~i3 & n285;
  assign n287 = ~i10 & n286;
  assign n288 = ~i7 & n287;
  assign n289 = n284 & ~n288;
  assign n290 = i10 & n286;
  assign n291 = n289 & ~n290;
  assign n292 = i2 & ~i11;
  assign n293 = n291 & ~n292;
  assign n294 = i2 & i11;
  assign n295 = ~i9 & n294;
  assign n296 = n293 & ~n295;
  assign n297 = i9 & n294;
  assign n298 = i0 & n297;
  assign n299 = n296 & ~n298;
  assign n300 = ~n155 & n299;
  assign n301 = ~n160 & ~n300;
  assign n302 = ~n166 & n301;
  assign n303 = ~n171 & n302;
  assign n304 = ~n179 & n303;
  assign n305 = ~n98 & ~n304;
  assign n306 = ~n183 & ~n305;
  assign n307 = ~n191 & n306;
  assign n308 = ~n197 & n307;
  assign n309 = ~n203 & n308;
  assign n310 = ~n207 & ~n309;
  assign n311 = ~n210 & ~n310;
  assign n312 = ~n220 & n311;
  assign n313 = ~n228 & n312;
  assign n314 = ~n235 & n313;
  assign n315 = ~n240 & n314;
  assign n316 = ~n245 & n315;
  assign n317 = ~n249 & n316;
  assign n318 = ~n253 & ~n317;
  assign n319 = ~n261 & ~n318;
  assign n320 = ~n265 & n319;
  assign i8 = ~n272 & n320;
endmodule


