// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 15:53:45 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8;
  wire n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
    n24, n25, n26;
  assign n10 = ~i0 & i3;
  assign n11 = i4 & n10;
  assign n12 = i5 & n11;
  assign n13 = i6 & n12;
  assign n14 = i3 & i4;
  assign n15 = i5 & n14;
  assign n16 = i6 & n15;
  assign n17 = ~i3 & ~i7;
  assign n18 = ~i4 & n17;
  assign n19 = i4 & n17;
  assign n20 = ~i6 & n19;
  assign n21 = ~n18 & ~n20;
  assign n22 = i6 & n19;
  assign n23 = ~i5 & n22;
  assign n24 = n21 & ~n23;
  assign n25 = ~i7 & n24;
  assign n26 = ~n13 & ~n25;
  assign i8 = ~n16 & n26;
endmodule


