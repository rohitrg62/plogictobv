// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:28:29 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8, i9, i10, i11  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8, i9, i10, i11;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
    n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
    n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n54, n55,
    n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
    n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
    n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
    n110, n111, n112, n113, n114, n115, n116, n117, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295;
  assign n13 = i0 & i1;
  assign n14 = i2 & n13;
  assign n15 = i3 & n14;
  assign n16 = i4 & n15;
  assign n17 = i5 & n16;
  assign n18 = ~i7 & n17;
  assign n19 = i1 & i2;
  assign n20 = i3 & n19;
  assign n21 = i4 & n20;
  assign n22 = i5 & n21;
  assign n23 = i7 & n22;
  assign n24 = i0 & i2;
  assign n25 = i3 & n24;
  assign n26 = i4 & n25;
  assign n27 = i5 & n26;
  assign n28 = i7 & n27;
  assign n29 = ~i4 & n15;
  assign n30 = i5 & n29;
  assign n31 = i7 & n30;
  assign n32 = ~i5 & ~i6;
  assign n33 = i5 & ~i6;
  assign n34 = ~i0 & n33;
  assign n35 = ~n32 & ~n34;
  assign n36 = i0 & n33;
  assign n37 = n35 & ~n36;
  assign n38 = ~i4 & i6;
  assign n39 = ~i5 & n38;
  assign n40 = n37 & ~n39;
  assign n41 = i5 & n38;
  assign n42 = n40 & ~n41;
  assign n43 = i4 & i6;
  assign n44 = ~i3 & n43;
  assign n45 = ~i5 & n44;
  assign n46 = ~i2 & n45;
  assign n47 = n42 & ~n46;
  assign n48 = i5 & n44;
  assign n49 = n47 & ~n48;
  assign n50 = ~n18 & n49;
  assign n51 = ~n23 & ~n50;
  assign n52 = ~n28 & n51;
  assign i11 = ~n31 & n52;
  assign n54 = ~i3 & n19;
  assign n55 = ~i4 & n54;
  assign n56 = ~i5 & n55;
  assign n57 = i6 & n56;
  assign n58 = i7 & n57;
  assign n59 = ~i0 & i1;
  assign n60 = i2 & n59;
  assign n61 = i3 & n60;
  assign n62 = i4 & n61;
  assign n63 = ~i5 & n62;
  assign n64 = i7 & n63;
  assign n65 = i0 & ~i1;
  assign n66 = i2 & n65;
  assign n67 = i3 & n66;
  assign n68 = i4 & n67;
  assign n69 = ~i5 & n68;
  assign n70 = i7 & n69;
  assign n71 = ~i3 & n14;
  assign n72 = i4 & n71;
  assign n73 = ~i5 & n72;
  assign n74 = ~i6 & n73;
  assign n75 = i7 & n74;
  assign n76 = i11 & n75;
  assign n77 = ~i7 & n27;
  assign n78 = i11 & n77;
  assign n79 = ~i0 & ~i1;
  assign n80 = i2 & n79;
  assign n81 = ~i4 & n80;
  assign n82 = ~i5 & n81;
  assign n83 = ~i6 & n82;
  assign n84 = i7 & n83;
  assign n85 = ~i4 & n25;
  assign n86 = i5 & n85;
  assign n87 = i2 & ~i3;
  assign n88 = ~i4 & n87;
  assign n89 = ~i5 & n88;
  assign n90 = ~i6 & n89;
  assign n91 = i7 & n90;
  assign n92 = i5 & n72;
  assign n93 = i7 & n92;
  assign n94 = i11 & n93;
  assign n95 = ~i2 & i11;
  assign n96 = i11 & ~n95;
  assign n97 = i2 & i11;
  assign n98 = ~i7 & n97;
  assign n99 = ~i5 & n98;
  assign n100 = n96 & ~n99;
  assign n101 = i5 & n98;
  assign n102 = n100 & ~n101;
  assign n103 = i7 & n97;
  assign n104 = i1 & n103;
  assign n105 = ~i5 & n104;
  assign n106 = n102 & ~n105;
  assign n107 = i5 & n104;
  assign n108 = n106 & ~n107;
  assign n109 = ~n58 & ~n108;
  assign n110 = ~n64 & n109;
  assign n111 = ~n17 & n110;
  assign n112 = ~n70 & n111;
  assign n113 = ~n76 & n112;
  assign n114 = ~n78 & n113;
  assign n115 = ~n84 & ~n114;
  assign n116 = ~n86 & n115;
  assign n117 = ~n91 & n116;
  assign i10 = ~n94 & ~n117;
  assign n119 = ~i3 & n13;
  assign n120 = i4 & n119;
  assign n121 = ~i5 & n120;
  assign n122 = i6 & n121;
  assign n123 = i7 & n122;
  assign n124 = i10 & n123;
  assign n125 = i11 & n124;
  assign n126 = i1 & ~i2;
  assign n127 = i3 & n126;
  assign n128 = ~i4 & n127;
  assign n129 = ~i5 & n128;
  assign n130 = i6 & n129;
  assign n131 = i7 & n130;
  assign n132 = i10 & n131;
  assign n133 = i2 & i3;
  assign n134 = i4 & n133;
  assign n135 = i5 & n134;
  assign n136 = ~i7 & n135;
  assign n137 = i10 & n136;
  assign n138 = ~i11 & n137;
  assign n139 = i7 & n73;
  assign n140 = i10 & n139;
  assign n141 = ~i0 & i2;
  assign n142 = i3 & n141;
  assign n143 = i4 & n142;
  assign n144 = ~i5 & n143;
  assign n145 = i7 & n144;
  assign n146 = i10 & n145;
  assign n147 = i0 & ~i2;
  assign n148 = i3 & n147;
  assign n149 = ~i4 & n148;
  assign n150 = ~i5 & n149;
  assign n151 = i6 & n150;
  assign n152 = i7 & n151;
  assign n153 = i10 & n152;
  assign n154 = n27 & ~i10;
  assign n155 = n27 & i10;
  assign n156 = ~i3 & n24;
  assign n157 = i4 & n156;
  assign n158 = ~i5 & n157;
  assign n159 = ~i10 & n158;
  assign n160 = i7 & n135;
  assign n161 = ~i10 & n160;
  assign n162 = i11 & n161;
  assign n163 = ~i4 & n133;
  assign n164 = i5 & n163;
  assign n165 = i7 & n164;
  assign n166 = i11 & n165;
  assign n167 = ~i4 & n14;
  assign n168 = i5 & n167;
  assign n169 = ~i11 & n168;
  assign n170 = ~i4 & n156;
  assign n171 = i5 & n170;
  assign n172 = i6 & n171;
  assign n173 = i7 & n172;
  assign n174 = ~i10 & n173;
  assign n175 = i11 & n174;
  assign n176 = i7 & n171;
  assign n177 = ~i10 & n176;
  assign n178 = i11 & n177;
  assign n179 = ~n125 & ~n132;
  assign n180 = ~n138 & n179;
  assign n181 = ~n140 & n180;
  assign n182 = ~n146 & n181;
  assign n183 = ~n153 & n182;
  assign n184 = ~n154 & ~n183;
  assign n185 = ~n155 & ~n184;
  assign n186 = ~n159 & ~n185;
  assign n187 = ~n154 & n186;
  assign n188 = ~n162 & ~n187;
  assign n189 = ~n166 & n188;
  assign n190 = ~n154 & ~n189;
  assign n191 = ~n169 & n190;
  assign n192 = ~n175 & ~n191;
  assign i9 = ~n178 & n192;
  assign n194 = i2 & i4;
  assign n195 = i5 & n194;
  assign n196 = ~i7 & n195;
  assign n197 = ~i9 & n196;
  assign n198 = ~i11 & n197;
  assign n199 = i0 & i3;
  assign n200 = i4 & n199;
  assign n201 = i5 & n200;
  assign n202 = i6 & n201;
  assign n203 = i7 & n202;
  assign n204 = i9 & n203;
  assign n205 = i10 & n204;
  assign n206 = ~i11 & n205;
  assign n207 = ~i6 & n195;
  assign n208 = ~i7 & n207;
  assign n209 = ~i10 & n208;
  assign n210 = i11 & n209;
  assign n211 = ~i9 & n207;
  assign n212 = ~i10 & n211;
  assign n213 = i11 & n212;
  assign n214 = i4 & n87;
  assign n215 = i5 & n214;
  assign n216 = i6 & n215;
  assign n217 = i7 & n216;
  assign n218 = i9 & n217;
  assign n219 = ~i10 & n218;
  assign n220 = i11 & n219;
  assign n221 = i0 & ~i3;
  assign n222 = i4 & n221;
  assign n223 = i5 & n222;
  assign n224 = i6 & n223;
  assign n225 = i7 & n224;
  assign n226 = i9 & n225;
  assign n227 = i10 & n226;
  assign n228 = i11 & n227;
  assign n229 = i6 & n195;
  assign n230 = i9 & n229;
  assign n231 = ~i10 & n230;
  assign n232 = ~i11 & n231;
  assign n233 = i3 & ~i4;
  assign n234 = i5 & n233;
  assign n235 = i6 & n234;
  assign n236 = i7 & n235;
  assign n237 = i9 & n236;
  assign n238 = i10 & n237;
  assign n239 = i11 & n238;
  assign n240 = i2 & ~i4;
  assign n241 = i5 & n240;
  assign n242 = i7 & n241;
  assign n243 = ~i9 & n242;
  assign n244 = i10 & n243;
  assign n245 = ~i10 & n207;
  assign n246 = ~i11 & n245;
  assign n247 = i7 & n207;
  assign n248 = ~i9 & n247;
  assign n249 = i10 & n248;
  assign n250 = ~i11 & n249;
  assign n251 = i5 & n88;
  assign n252 = ~i6 & n251;
  assign n253 = i7 & n252;
  assign n254 = i9 & n253;
  assign n255 = ~i10 & n254;
  assign n256 = i11 & n255;
  assign n257 = i6 & n241;
  assign n258 = i7 & n257;
  assign n259 = i9 & n258;
  assign n260 = i10 & n259;
  assign n261 = ~i11 & n260;
  assign n262 = ~i6 & n241;
  assign n263 = i7 & n262;
  assign n264 = i10 & n263;
  assign n265 = ~i11 & n264;
  assign n266 = ~i9 & n252;
  assign n267 = ~i10 & n266;
  assign n268 = i5 & ~n33;
  assign n269 = i5 & i6;
  assign n270 = ~i2 & n269;
  assign n271 = n268 & ~n270;
  assign n272 = i2 & n269;
  assign n273 = ~i10 & n272;
  assign n274 = n271 & ~n273;
  assign n275 = i10 & n272;
  assign n276 = ~i4 & n275;
  assign n277 = ~i11 & n276;
  assign n278 = n274 & ~n277;
  assign n279 = i11 & n276;
  assign n280 = ~i9 & n279;
  assign n281 = n278 & ~n280;
  assign n282 = ~n198 & n281;
  assign n283 = ~n206 & ~n282;
  assign n284 = ~n210 & n283;
  assign n285 = ~n213 & n284;
  assign n286 = ~n220 & n285;
  assign n287 = ~n228 & n286;
  assign n288 = ~n232 & n287;
  assign n289 = ~n239 & n288;
  assign n290 = ~n244 & n289;
  assign n291 = ~n246 & ~n290;
  assign n292 = ~n250 & ~n291;
  assign n293 = ~n256 & n292;
  assign n294 = ~n261 & ~n293;
  assign n295 = ~n265 & ~n294;
  assign i8 = n267 | n295;
endmodule


