// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:27:54 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8, i9, i10, i11  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8, i9, i10, i11;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
    n27, n28, n29, n30, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
    n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
    n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291;
  assign n13 = i1 & ~i5;
  assign n14 = ~i0 & n13;
  assign n15 = i2 & n14;
  assign n16 = i6 & n15;
  assign n17 = i1 & ~n16;
  assign n18 = i0 & n13;
  assign n19 = ~i3 & n18;
  assign n20 = n17 & ~n19;
  assign n21 = i3 & n18;
  assign n22 = n20 & ~n21;
  assign n23 = i1 & i5;
  assign n24 = ~i2 & n23;
  assign n25 = n22 & ~n24;
  assign n26 = i2 & n23;
  assign n27 = ~i0 & n26;
  assign n28 = n25 & ~n27;
  assign n29 = i0 & n26;
  assign n30 = ~i3 & n29;
  assign i8 = ~n28 | n30;
  assign n32 = i2 & i3;
  assign n33 = ~i4 & n32;
  assign n34 = ~i5 & n33;
  assign n35 = i7 & n34;
  assign n36 = i7 & n33;
  assign n37 = ~i8 & n36;
  assign n38 = i1 & i2;
  assign n39 = i3 & n38;
  assign n40 = ~i4 & n39;
  assign n41 = i5 & n40;
  assign n42 = i7 & n41;
  assign n43 = i8 & n42;
  assign n44 = i0 & i2;
  assign n45 = i3 & n44;
  assign n46 = i4 & n45;
  assign n47 = ~i5 & n46;
  assign n48 = i7 & n47;
  assign n49 = i4 & n32;
  assign n50 = i5 & n49;
  assign n51 = ~i7 & n50;
  assign n52 = i8 & n51;
  assign n53 = i7 & n46;
  assign n54 = ~i8 & n53;
  assign n55 = i4 & n39;
  assign n56 = ~i5 & n55;
  assign n57 = i7 & n56;
  assign n58 = ~i8 & n57;
  assign n59 = i0 & i1;
  assign n60 = i2 & n59;
  assign n61 = i4 & n60;
  assign n62 = i5 & n61;
  assign n63 = ~i7 & n62;
  assign n64 = i8 & n63;
  assign n65 = ~i4 & n45;
  assign n66 = i5 & n65;
  assign n67 = i7 & n66;
  assign n68 = i8 & n67;
  assign n69 = ~n35 & ~n37;
  assign n70 = ~n43 & n69;
  assign n71 = ~n48 & n70;
  assign n72 = ~n52 & n71;
  assign n73 = ~n54 & n72;
  assign n74 = ~n58 & n73;
  assign n75 = ~n64 & n74;
  assign i11 = ~n68 & n75;
  assign n77 = n36 & i11;
  assign n78 = i4 & n44;
  assign n79 = ~i5 & n78;
  assign n80 = i7 & n79;
  assign n81 = ~i11 & n80;
  assign n82 = i7 & n78;
  assign n83 = ~i8 & n82;
  assign n84 = ~i11 & n83;
  assign n85 = i4 & n38;
  assign n86 = ~i5 & n85;
  assign n87 = i7 & n86;
  assign n88 = ~i8 & n87;
  assign n89 = ~i11 & n88;
  assign n90 = ~i7 & n78;
  assign n91 = ~i8 & n90;
  assign n92 = i11 & n91;
  assign n93 = i8 & n66;
  assign n94 = i4 & i5;
  assign n95 = ~i4 & ~i5;
  assign n96 = i4 & ~i5;
  assign n97 = ~i2 & n96;
  assign n98 = ~i11 & n97;
  assign n99 = ~n95 & ~n98;
  assign n100 = i11 & n97;
  assign n101 = ~i0 & n100;
  assign n102 = n99 & ~n101;
  assign n103 = i2 & n96;
  assign n104 = i7 & n103;
  assign n105 = i11 & n104;
  assign n106 = n102 & ~n105;
  assign n107 = ~i4 & i5;
  assign n108 = ~i8 & n107;
  assign n109 = n106 & ~n108;
  assign n110 = i8 & n107;
  assign n111 = ~i2 & n110;
  assign n112 = ~i1 & n111;
  assign n113 = ~i7 & n112;
  assign n114 = n109 & ~n113;
  assign n115 = i7 & n112;
  assign n116 = n114 & ~n115;
  assign n117 = i1 & n111;
  assign n118 = ~i6 & n117;
  assign n119 = n116 & ~n118;
  assign n120 = i2 & n110;
  assign n121 = ~i3 & n120;
  assign n122 = i7 & n121;
  assign n123 = n119 & ~n122;
  assign n124 = ~n94 & n123;
  assign n125 = ~n77 & n124;
  assign n126 = ~n81 & ~n125;
  assign n127 = ~n84 & n126;
  assign n128 = ~n89 & n127;
  assign n129 = ~n92 & n128;
  assign i10 = ~n93 & n129;
  assign n131 = i3 & ~i4;
  assign n132 = ~i5 & n131;
  assign n133 = ~i6 & n132;
  assign n134 = i7 & n133;
  assign n135 = i11 & n134;
  assign n136 = i2 & ~i4;
  assign n137 = ~i5 & n136;
  assign n138 = i6 & n137;
  assign n139 = ~i11 & n138;
  assign n140 = i6 & n136;
  assign n141 = ~i8 & n140;
  assign n142 = ~i11 & n141;
  assign n143 = i2 & i4;
  assign n144 = i6 & n143;
  assign n145 = i10 & n144;
  assign n146 = i11 & n145;
  assign n147 = i3 & ~i5;
  assign n148 = ~i6 & n147;
  assign n149 = i7 & n148;
  assign n150 = ~i10 & n149;
  assign n151 = i11 & n150;
  assign n152 = i3 & n59;
  assign n153 = ~i4 & n152;
  assign n154 = i5 & n153;
  assign n155 = i6 & n154;
  assign n156 = ~i7 & n155;
  assign n157 = i8 & n156;
  assign n158 = ~i10 & n157;
  assign n159 = ~i6 & n136;
  assign n160 = ~i10 & n159;
  assign n161 = ~i11 & n160;
  assign n162 = i2 & ~i5;
  assign n163 = i6 & n162;
  assign n164 = ~i10 & n163;
  assign n165 = ~i11 & n164;
  assign n166 = i3 & i4;
  assign n167 = ~i6 & n166;
  assign n168 = ~i7 & n167;
  assign n169 = i10 & n168;
  assign n170 = i11 & n169;
  assign n171 = i4 & n59;
  assign n172 = i5 & n171;
  assign n173 = ~i6 & n172;
  assign n174 = ~i7 & n173;
  assign n175 = i8 & n174;
  assign n176 = i10 & n175;
  assign n177 = i11 & n176;
  assign n178 = i5 & n152;
  assign n179 = ~i6 & n178;
  assign n180 = i7 & n179;
  assign n181 = i8 & n180;
  assign n182 = i11 & n181;
  assign n183 = i2 & ~i6;
  assign n184 = ~i7 & n183;
  assign n185 = ~i11 & n184;
  assign n186 = ~i8 & n183;
  assign n187 = ~i10 & n186;
  assign n188 = ~i11 & n187;
  assign n189 = ~i6 & n162;
  assign n190 = ~i10 & n189;
  assign n191 = ~i11 & n190;
  assign n192 = i2 & i6;
  assign n193 = ~i7 & n192;
  assign n194 = ~i11 & n193;
  assign n195 = i1 & i3;
  assign n196 = i4 & n195;
  assign n197 = ~i5 & n196;
  assign n198 = ~i6 & n197;
  assign n199 = i7 & n198;
  assign n200 = ~i8 & n199;
  assign n201 = i10 & n200;
  assign n202 = i11 & n201;
  assign n203 = i1 & i4;
  assign n204 = ~i5 & n203;
  assign n205 = ~i6 & n204;
  assign n206 = ~i7 & n205;
  assign n207 = ~i8 & n206;
  assign n208 = i10 & n207;
  assign n209 = i11 & n208;
  assign n210 = i8 & n179;
  assign n211 = i10 & n210;
  assign n212 = i11 & n211;
  assign n213 = i0 & i3;
  assign n214 = ~i4 & n213;
  assign n215 = i5 & n214;
  assign n216 = ~i6 & n215;
  assign n217 = i7 & n216;
  assign n218 = i8 & n217;
  assign n219 = i10 & n218;
  assign n220 = i11 & n219;
  assign n221 = ~i8 & n193;
  assign n222 = ~i10 & n221;
  assign n223 = ~i10 & n140;
  assign n224 = ~i11 & n223;
  assign n225 = ~i4 & n195;
  assign n226 = i5 & n225;
  assign n227 = ~i6 & n226;
  assign n228 = i7 & n227;
  assign n229 = i8 & n228;
  assign n230 = i10 & n229;
  assign n231 = i11 & n230;
  assign n232 = i3 & i5;
  assign n233 = ~i6 & n232;
  assign n234 = ~i7 & n233;
  assign n235 = i8 & n234;
  assign n236 = i10 & n235;
  assign n237 = i11 & n236;
  assign n238 = i0 & ~i4;
  assign n239 = i5 & n238;
  assign n240 = ~i6 & n239;
  assign n241 = ~i7 & n240;
  assign n242 = i8 & n241;
  assign n243 = i10 & n242;
  assign n244 = i11 & n243;
  assign n245 = i1 & ~i4;
  assign n246 = i5 & n245;
  assign n247 = ~i6 & n246;
  assign n248 = ~i7 & n247;
  assign n249 = i8 & n248;
  assign n250 = i10 & n249;
  assign n251 = i11 & n250;
  assign n252 = ~i11 & n183;
  assign n253 = i2 & ~n252;
  assign n254 = i11 & n183;
  assign n255 = ~i7 & n254;
  assign n256 = ~i10 & n255;
  assign n257 = n253 & ~n256;
  assign n258 = i10 & n255;
  assign n259 = ~i4 & n258;
  assign n260 = n257 & ~n259;
  assign n261 = i7 & n192;
  assign n262 = ~i11 & n261;
  assign n263 = ~i3 & n262;
  assign n264 = i5 & n263;
  assign n265 = n260 & ~n264;
  assign n266 = i11 & n261;
  assign n267 = n265 & ~n266;
  assign n268 = ~n135 & ~n267;
  assign n269 = ~n139 & n268;
  assign n270 = ~n142 & n269;
  assign n271 = ~n146 & ~n270;
  assign n272 = ~n151 & ~n271;
  assign n273 = ~n158 & n272;
  assign n274 = ~n161 & ~n273;
  assign n275 = ~n165 & ~n274;
  assign n276 = ~n170 & n275;
  assign n277 = ~n177 & n276;
  assign n278 = ~n182 & n277;
  assign n279 = ~n185 & ~n278;
  assign n280 = ~n188 & n279;
  assign n281 = ~n191 & n280;
  assign n282 = ~n194 & ~n281;
  assign n283 = ~n202 & n282;
  assign n284 = ~n209 & n283;
  assign n285 = ~n212 & n284;
  assign n286 = ~n220 & n285;
  assign n287 = ~n222 & n286;
  assign n288 = ~n224 & n287;
  assign n289 = ~n231 & n288;
  assign n290 = ~n237 & n289;
  assign n291 = ~n244 & n290;
  assign i9 = ~n251 & n291;
endmodule


