// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:27:10 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8, i9, i10, i11  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8, i9, i10, i11;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
    n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
    n41, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
    n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
    n84, n85, n86, n87, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276;
  assign n13 = ~i0 & ~i1;
  assign n14 = i2 & n13;
  assign n15 = ~i3 & n14;
  assign n16 = i6 & n15;
  assign n17 = i1 & ~i4;
  assign n18 = ~i5 & n17;
  assign n19 = i6 & n18;
  assign n20 = ~i7 & n19;
  assign n21 = i3 & n13;
  assign n22 = i6 & n21;
  assign n23 = ~i7 & n22;
  assign n24 = i0 & ~i1;
  assign n25 = ~i4 & n24;
  assign n26 = i6 & n25;
  assign n27 = ~i7 & n26;
  assign n28 = ~i1 & ~i4;
  assign n29 = ~i2 & n28;
  assign n30 = ~i3 & n29;
  assign n31 = ~n17 & ~n30;
  assign n32 = ~i3 & i4;
  assign n33 = n31 & ~n32;
  assign n34 = i3 & i4;
  assign n35 = ~i2 & n34;
  assign n36 = n33 & ~n35;
  assign n37 = i2 & n34;
  assign n38 = n36 & ~n37;
  assign n39 = ~n16 & n38;
  assign n40 = ~n20 & ~n39;
  assign n41 = ~n23 & n40;
  assign i11 = ~n27 & n41;
  assign n43 = ~i0 & i1;
  assign n44 = ~i3 & n43;
  assign n45 = ~i4 & n44;
  assign n46 = ~i5 & n45;
  assign n47 = i6 & n46;
  assign n48 = i11 & n47;
  assign n49 = i0 & i1;
  assign n50 = ~i3 & n49;
  assign n51 = ~i4 & n50;
  assign n52 = ~i5 & n51;
  assign n53 = i6 & n52;
  assign n54 = i11 & n53;
  assign n55 = ~i5 & n50;
  assign n56 = i6 & n55;
  assign n57 = ~i7 & n56;
  assign n58 = i11 & n57;
  assign n59 = i6 & n44;
  assign n60 = ~i7 & n59;
  assign n61 = i6 & n51;
  assign n62 = ~i7 & n61;
  assign n63 = ~i11 & n62;
  assign n64 = ~i1 & ~i11;
  assign n65 = ~i1 & i11;
  assign n66 = ~i0 & n65;
  assign n67 = ~n64 & ~n66;
  assign n68 = i0 & n65;
  assign n69 = ~i2 & n68;
  assign n70 = n67 & ~n69;
  assign n71 = i2 & n68;
  assign n72 = ~i6 & n71;
  assign n73 = i4 & n72;
  assign n74 = n70 & ~n73;
  assign n75 = i1 & ~i3;
  assign n76 = ~i5 & n75;
  assign n77 = n74 & ~n76;
  assign n78 = i1 & i3;
  assign n79 = ~i11 & n78;
  assign n80 = ~i6 & n79;
  assign n81 = n77 & ~n80;
  assign n82 = i11 & n78;
  assign n83 = n81 & ~n82;
  assign n84 = ~n48 & ~n83;
  assign n85 = ~n54 & n84;
  assign n86 = ~n58 & n85;
  assign n87 = ~n60 & n86;
  assign i9 = ~n63 & n87;
  assign n89 = i2 & n43;
  assign n90 = i3 & n89;
  assign n91 = ~i5 & n90;
  assign n92 = i6 & n91;
  assign n93 = ~i7 & n92;
  assign n94 = i9 & n93;
  assign n95 = i11 & n94;
  assign n96 = ~i2 & n49;
  assign n97 = ~i3 & n96;
  assign n98 = ~i5 & n97;
  assign n99 = i6 & n98;
  assign n100 = ~i7 & n99;
  assign n101 = ~i9 & n100;
  assign n102 = i11 & n101;
  assign n103 = i2 & n49;
  assign n104 = ~i3 & n103;
  assign n105 = ~i5 & n104;
  assign n106 = i6 & n105;
  assign n107 = ~i7 & n106;
  assign n108 = ~i9 & n107;
  assign n109 = i11 & n108;
  assign n110 = ~i2 & n43;
  assign n111 = i3 & n110;
  assign n112 = ~i4 & n111;
  assign n113 = i6 & n112;
  assign n114 = ~i7 & n113;
  assign n115 = i9 & n114;
  assign n116 = i11 & n115;
  assign n117 = ~i4 & n90;
  assign n118 = i6 & n117;
  assign n119 = ~i7 & n118;
  assign n120 = i9 & n119;
  assign n121 = i11 & n120;
  assign n122 = ~i5 & n111;
  assign n123 = i6 & n122;
  assign n124 = ~i7 & n123;
  assign n125 = i9 & n124;
  assign n126 = i11 & n125;
  assign n127 = ~i4 & n97;
  assign n128 = i6 & n127;
  assign n129 = ~i7 & n128;
  assign n130 = ~i9 & n129;
  assign n131 = i11 & n130;
  assign n132 = i1 & ~i2;
  assign n133 = i1 & ~n132;
  assign n134 = i1 & i2;
  assign n135 = ~i11 & n134;
  assign n136 = i6 & n135;
  assign n137 = n133 & ~n136;
  assign n138 = i11 & n134;
  assign n139 = i5 & n138;
  assign n140 = ~i6 & n139;
  assign n141 = n137 & ~n140;
  assign n142 = i6 & n139;
  assign n143 = ~i9 & n142;
  assign n144 = ~i0 & n143;
  assign n145 = i3 & n144;
  assign n146 = n141 & ~n145;
  assign n147 = i0 & n143;
  assign n148 = n146 & ~n147;
  assign n149 = ~n95 & n148;
  assign n150 = ~n102 & ~n149;
  assign n151 = ~n109 & ~n150;
  assign n152 = ~n116 & ~n151;
  assign n153 = ~n121 & ~n152;
  assign n154 = ~n126 & ~n153;
  assign i10 = ~n131 & n154;
  assign n156 = i2 & n24;
  assign n157 = ~i3 & n156;
  assign n158 = ~i6 & n157;
  assign n159 = ~i7 & n158;
  assign n160 = i9 & n159;
  assign n161 = i11 & n160;
  assign n162 = i3 & n156;
  assign n163 = ~i6 & n162;
  assign n164 = ~i7 & n163;
  assign n165 = i9 & n164;
  assign n166 = i11 & n165;
  assign n167 = i6 & n97;
  assign n168 = ~i9 & n167;
  assign n169 = i10 & n168;
  assign n170 = i11 & n169;
  assign n171 = ~i5 & n112;
  assign n172 = ~i7 & n171;
  assign n173 = i9 & n172;
  assign n174 = i10 & n173;
  assign n175 = i11 & n174;
  assign n176 = ~i5 & n49;
  assign n177 = i6 & n176;
  assign n178 = ~i7 & n177;
  assign n179 = i11 & n178;
  assign n180 = ~i2 & n24;
  assign n181 = i3 & n180;
  assign n182 = i6 & n181;
  assign n183 = i9 & n182;
  assign n184 = ~i11 & n183;
  assign n185 = ~i3 & n24;
  assign n186 = ~i4 & n185;
  assign n187 = i6 & n186;
  assign n188 = i11 & n187;
  assign n189 = i6 & n104;
  assign n190 = ~i9 & n189;
  assign n191 = ~i10 & n190;
  assign n192 = i11 & n191;
  assign n193 = i3 & n14;
  assign n194 = ~i6 & n193;
  assign n195 = ~i7 & n194;
  assign n196 = i11 & n195;
  assign n197 = ~i5 & n117;
  assign n198 = ~i6 & n197;
  assign n199 = ~i7 & n198;
  assign n200 = i9 & n199;
  assign n201 = ~i10 & n200;
  assign n202 = i11 & n201;
  assign n203 = ~i2 & n13;
  assign n204 = i3 & n203;
  assign n205 = ~i7 & n204;
  assign n206 = i11 & n205;
  assign n207 = ~i7 & n98;
  assign n208 = i9 & n207;
  assign n209 = i10 & n208;
  assign n210 = i11 & n209;
  assign n211 = ~i5 & n43;
  assign n212 = i6 & n211;
  assign n213 = ~i7 & n212;
  assign n214 = i11 & n213;
  assign n215 = i6 & n185;
  assign n216 = ~i7 & n215;
  assign n217 = ~i5 & n44;
  assign n218 = i6 & n217;
  assign n219 = i9 & n218;
  assign n220 = i11 & n219;
  assign n221 = i6 & n193;
  assign n222 = i11 & n221;
  assign n223 = i0 & ~i4;
  assign n224 = i6 & n223;
  assign n225 = ~i7 & n224;
  assign n226 = i11 & n225;
  assign n227 = i3 & n24;
  assign n228 = i6 & n227;
  assign n229 = ~i7 & n228;
  assign n230 = i11 & n229;
  assign n231 = i6 & n204;
  assign n232 = ~i11 & n231;
  assign n233 = i6 & n14;
  assign n234 = ~i11 & n233;
  assign n235 = i6 & n162;
  assign n236 = i9 & n235;
  assign n237 = ~i11 & n236;
  assign n238 = ~i4 & ~i7;
  assign n239 = ~i11 & n238;
  assign n240 = ~i0 & n239;
  assign n241 = ~i1 & n240;
  assign n242 = i11 & n238;
  assign n243 = i0 & n242;
  assign n244 = ~n241 & ~n243;
  assign n245 = i4 & ~i7;
  assign n246 = ~i10 & n245;
  assign n247 = n244 & ~n246;
  assign n248 = i10 & n245;
  assign n249 = i5 & n248;
  assign n250 = n247 & ~n249;
  assign n251 = ~i3 & i7;
  assign n252 = i11 & n251;
  assign n253 = n250 & ~n252;
  assign n254 = i3 & i7;
  assign n255 = n253 & ~n254;
  assign n256 = ~n161 & ~n255;
  assign n257 = ~n166 & ~n256;
  assign n258 = ~n170 & ~n257;
  assign n259 = ~n175 & ~n258;
  assign n260 = ~n179 & n259;
  assign n261 = ~n184 & ~n260;
  assign n262 = ~n188 & n261;
  assign n263 = ~n192 & n262;
  assign n264 = ~n196 & n263;
  assign n265 = ~n202 & ~n264;
  assign n266 = ~n206 & n265;
  assign n267 = ~n210 & n266;
  assign n268 = ~n214 & ~n267;
  assign n269 = ~n216 & n268;
  assign n270 = ~n220 & n269;
  assign n271 = ~n179 & ~n270;
  assign n272 = ~n222 & ~n271;
  assign n273 = ~n226 & ~n272;
  assign n274 = ~n230 & n273;
  assign n275 = ~n232 & n274;
  assign n276 = ~n234 & n275;
  assign i8 = ~n237 & ~n276;
endmodule


