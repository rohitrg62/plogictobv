// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:27:09 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8, i9, i10, i11  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8, i9, i10, i11;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
    n27, n28, n29, n30, n31, n32, n34, n35, n36, n37, n38, n39, n40, n41,
    n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
    n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333;
  assign n13 = ~i0 & ~i1;
  assign n14 = i2 & n13;
  assign n15 = ~i3 & n14;
  assign n16 = ~i4 & n15;
  assign n17 = ~i5 & n16;
  assign n18 = ~i6 & n17;
  assign n19 = ~i7 & n18;
  assign n20 = ~i1 & ~i5;
  assign n21 = ~i4 & n20;
  assign n22 = ~i0 & n21;
  assign n23 = ~i7 & n22;
  assign n24 = ~i3 & n23;
  assign n25 = i7 & n22;
  assign n26 = ~n24 & ~n25;
  assign n27 = i4 & n20;
  assign n28 = n26 & ~n27;
  assign n29 = ~i1 & i5;
  assign n30 = n28 & ~n29;
  assign n31 = i1 & i5;
  assign n32 = n30 & ~n31;
  assign i8 = ~n19 & ~n32;
  assign n34 = ~i2 & n13;
  assign n35 = i3 & n34;
  assign n36 = ~i4 & n35;
  assign n37 = ~i5 & n36;
  assign n38 = ~i6 & n37;
  assign n39 = i3 & n13;
  assign n40 = ~i4 & n39;
  assign n41 = ~i5 & n40;
  assign n42 = ~i6 & n41;
  assign n43 = ~i8 & n42;
  assign n44 = i3 & n14;
  assign n45 = ~i4 & n44;
  assign n46 = ~i5 & n45;
  assign n47 = i6 & n46;
  assign n48 = i8 & n47;
  assign n49 = ~i0 & n20;
  assign n50 = ~i3 & n49;
  assign n51 = i3 & n49;
  assign n52 = ~n50 & ~n51;
  assign n53 = i0 & n20;
  assign n54 = ~i7 & n53;
  assign n55 = i4 & n54;
  assign n56 = i3 & n55;
  assign n57 = n52 & ~n56;
  assign n58 = i7 & n53;
  assign n59 = ~i3 & n58;
  assign n60 = n57 & ~n59;
  assign n61 = i3 & n58;
  assign n62 = ~i4 & n61;
  assign n63 = n60 & ~n62;
  assign n64 = ~n29 & n63;
  assign n65 = i1 & ~i4;
  assign n66 = i0 & n65;
  assign n67 = i8 & n66;
  assign n68 = n64 & ~n67;
  assign n69 = i1 & i4;
  assign n70 = ~i5 & n69;
  assign n71 = n68 & ~n70;
  assign n72 = i5 & n69;
  assign n73 = ~i0 & n72;
  assign n74 = n71 & ~n73;
  assign n75 = ~n38 & ~n74;
  assign n76 = ~n43 & n75;
  assign i9 = ~n48 & n76;
  assign n78 = i1 & i2;
  assign n79 = ~i3 & n78;
  assign n80 = i6 & n79;
  assign n81 = i7 & n80;
  assign n82 = i8 & n81;
  assign n83 = i9 & n82;
  assign n84 = ~i0 & i1;
  assign n85 = i2 & n84;
  assign n86 = ~i3 & n85;
  assign n87 = i6 & n86;
  assign n88 = i8 & n87;
  assign n89 = i1 & ~i2;
  assign n90 = ~i3 & n89;
  assign n91 = ~i6 & n90;
  assign n92 = i7 & n91;
  assign n93 = i9 & n92;
  assign n94 = ~i2 & n84;
  assign n95 = ~i3 & n94;
  assign n96 = ~i6 & n95;
  assign n97 = ~i9 & n96;
  assign n98 = i3 & n85;
  assign n99 = ~i6 & n98;
  assign n100 = ~i7 & n99;
  assign n101 = i8 & n100;
  assign n102 = ~i9 & n101;
  assign n103 = i0 & i1;
  assign n104 = i2 & n103;
  assign n105 = ~i3 & n104;
  assign n106 = ~i6 & n105;
  assign n107 = i7 & n106;
  assign n108 = i8 & n107;
  assign n109 = ~i9 & n108;
  assign n110 = ~i7 & n91;
  assign n111 = ~i9 & n110;
  assign n112 = ~i2 & n103;
  assign n113 = ~i3 & n112;
  assign n114 = i6 & n113;
  assign n115 = i7 & n114;
  assign n116 = ~i8 & n115;
  assign n117 = ~i9 & n116;
  assign n118 = ~i7 & n114;
  assign n119 = i8 & n118;
  assign n120 = i9 & n119;
  assign n121 = ~i6 & n94;
  assign n122 = ~i8 & n121;
  assign n123 = ~i9 & n122;
  assign n124 = i1 & i3;
  assign n125 = i6 & n124;
  assign n126 = ~i8 & n125;
  assign n127 = i9 & n126;
  assign n128 = ~i3 & n84;
  assign n129 = ~i6 & n128;
  assign n130 = ~i8 & n129;
  assign n131 = ~i7 & n106;
  assign n132 = i8 & n131;
  assign n133 = i9 & n132;
  assign n134 = i6 & n98;
  assign n135 = i7 & n134;
  assign n136 = i8 & n135;
  assign n137 = ~i9 & n136;
  assign n138 = i3 & n112;
  assign n139 = ~i6 & n138;
  assign n140 = ~i7 & n139;
  assign n141 = i8 & n140;
  assign n142 = ~i9 & n141;
  assign n143 = i3 & n94;
  assign n144 = i6 & n143;
  assign n145 = i7 & n144;
  assign n146 = i8 & n145;
  assign n147 = i9 & n146;
  assign n148 = ~i6 & n84;
  assign n149 = ~i8 & n148;
  assign n150 = ~i9 & n149;
  assign n151 = i7 & n99;
  assign n152 = i8 & n151;
  assign n153 = i9 & n152;
  assign n154 = ~i6 & n143;
  assign n155 = i7 & n154;
  assign n156 = i8 & n155;
  assign n157 = ~i9 & n156;
  assign n158 = ~i7 & n144;
  assign n159 = i8 & n158;
  assign n160 = ~i9 & n159;
  assign n161 = ~i6 & n89;
  assign n162 = ~i7 & n161;
  assign n163 = ~i8 & n162;
  assign n164 = ~i9 & n163;
  assign n165 = ~i3 & n103;
  assign n166 = i6 & n165;
  assign n167 = i7 & n166;
  assign n168 = ~i8 & n167;
  assign n169 = ~i9 & n168;
  assign n170 = i3 & n89;
  assign n171 = ~i6 & n170;
  assign n172 = i7 & n171;
  assign n173 = i8 & n172;
  assign n174 = ~i9 & n173;
  assign n175 = i1 & ~i3;
  assign n176 = ~i6 & n175;
  assign n177 = ~i8 & n176;
  assign n178 = i9 & n177;
  assign n179 = i3 & n78;
  assign n180 = i6 & n179;
  assign n181 = i7 & n180;
  assign n182 = i8 & n181;
  assign n183 = ~i9 & n182;
  assign n184 = ~i7 & n154;
  assign n185 = i8 & n184;
  assign n186 = i9 & n185;
  assign n187 = ~i9 & n115;
  assign n188 = ~i7 & n80;
  assign n189 = i8 & n188;
  assign n190 = ~i9 & n189;
  assign n191 = i8 & n139;
  assign n192 = i9 & n191;
  assign n193 = i3 & n104;
  assign n194 = i6 & n193;
  assign n195 = ~i7 & n194;
  assign n196 = i8 & n195;
  assign n197 = ~i9 & n196;
  assign n198 = i8 & n194;
  assign n199 = i9 & n198;
  assign n200 = i6 & n112;
  assign n201 = i7 & n200;
  assign n202 = ~i8 & n201;
  assign n203 = ~i9 & n202;
  assign n204 = i6 & n103;
  assign n205 = i7 & n204;
  assign n206 = ~i8 & n205;
  assign n207 = ~i9 & n206;
  assign n208 = ~i7 & n176;
  assign n209 = ~i8 & n208;
  assign n210 = ~i9 & n209;
  assign n211 = i1 & ~i6;
  assign n212 = ~i7 & n211;
  assign n213 = ~i8 & n212;
  assign n214 = ~i9 & n213;
  assign n215 = ~i7 & n134;
  assign n216 = i8 & n215;
  assign n217 = i9 & n216;
  assign n218 = ~n83 & ~n88;
  assign n219 = ~n93 & n218;
  assign n220 = ~n97 & n219;
  assign n221 = ~n96 & n220;
  assign n222 = ~n102 & n221;
  assign n223 = ~n109 & n222;
  assign n224 = ~n111 & n223;
  assign n225 = ~n117 & n224;
  assign n226 = ~n120 & n225;
  assign n227 = ~n123 & n226;
  assign n228 = ~n127 & n227;
  assign n229 = ~n130 & n228;
  assign n230 = ~n133 & n229;
  assign n231 = ~n137 & n230;
  assign n232 = ~n142 & n231;
  assign n233 = ~n147 & n232;
  assign n234 = ~n150 & n233;
  assign n235 = ~n153 & n234;
  assign n236 = ~n157 & n235;
  assign n237 = ~n160 & n236;
  assign n238 = ~n164 & n237;
  assign n239 = ~n169 & n238;
  assign n240 = ~n174 & n239;
  assign n241 = ~n178 & n240;
  assign n242 = ~n183 & n241;
  assign n243 = ~n186 & n242;
  assign n244 = ~n187 & n243;
  assign n245 = ~n190 & n244;
  assign n246 = ~n192 & n245;
  assign n247 = ~n197 & n246;
  assign n248 = ~n199 & n247;
  assign n249 = ~n203 & n248;
  assign n250 = ~n207 & n249;
  assign n251 = ~n210 & n250;
  assign n252 = ~n214 & n251;
  assign i10 = ~n217 & n252;
  assign n254 = i0 & ~i1;
  assign n255 = ~i2 & n254;
  assign n256 = ~i3 & n255;
  assign n257 = ~i5 & n256;
  assign n258 = ~i6 & n257;
  assign n259 = i3 & n254;
  assign n260 = ~i5 & n259;
  assign n261 = i6 & n260;
  assign n262 = ~i8 & n261;
  assign n263 = i9 & n262;
  assign n264 = i7 & n165;
  assign n265 = ~i8 & n264;
  assign n266 = i9 & n265;
  assign n267 = i3 & n255;
  assign n268 = ~i5 & n267;
  assign n269 = ~i6 & n268;
  assign n270 = ~i8 & n269;
  assign n271 = i9 & n270;
  assign n272 = i2 & n254;
  assign n273 = ~i3 & n272;
  assign n274 = ~i5 & n273;
  assign n275 = i6 & n274;
  assign n276 = i8 & n275;
  assign n277 = ~i6 & n260;
  assign n278 = ~i8 & n277;
  assign n279 = i9 & n278;
  assign n280 = i8 & n269;
  assign n281 = i9 & n280;
  assign n282 = i3 & n272;
  assign n283 = ~i5 & n282;
  assign n284 = i6 & n283;
  assign n285 = i8 & n284;
  assign n286 = i9 & n285;
  assign n287 = ~i5 & n272;
  assign n288 = i6 & n287;
  assign n289 = i8 & n288;
  assign n290 = ~i9 & n289;
  assign n291 = ~i7 & n165;
  assign n292 = ~i8 & n291;
  assign n293 = i9 & n292;
  assign n294 = ~i5 & n255;
  assign n295 = ~i6 & n294;
  assign n296 = ~i9 & n295;
  assign n297 = ~i6 & n254;
  assign n298 = i8 & n297;
  assign n299 = ~n13 & ~n298;
  assign n300 = i6 & n254;
  assign n301 = ~i3 & n300;
  assign n302 = i10 & n301;
  assign n303 = n299 & ~n302;
  assign n304 = i3 & n300;
  assign n305 = n303 & ~n304;
  assign n306 = i1 & ~i7;
  assign n307 = i3 & n306;
  assign n308 = ~i5 & n307;
  assign n309 = i4 & n308;
  assign n310 = i0 & n309;
  assign n311 = n305 & ~n310;
  assign n312 = i5 & n307;
  assign n313 = n311 & ~n312;
  assign n314 = i1 & i7;
  assign n315 = ~i3 & n314;
  assign n316 = n313 & ~n315;
  assign n317 = i3 & n314;
  assign n318 = ~i8 & n317;
  assign n319 = ~i9 & n318;
  assign n320 = n316 & ~n319;
  assign n321 = i9 & n318;
  assign n322 = ~i0 & n321;
  assign n323 = n320 & ~n322;
  assign n324 = ~n258 & ~n323;
  assign n325 = ~n263 & n324;
  assign n326 = ~n266 & n325;
  assign n327 = ~n271 & ~n326;
  assign n328 = ~n276 & ~n327;
  assign n329 = ~n279 & ~n328;
  assign n330 = ~n281 & ~n329;
  assign n331 = ~n286 & n330;
  assign n332 = ~n290 & n331;
  assign n333 = ~n293 & ~n332;
  assign i11 = ~n296 & ~n333;
endmodule


