// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 15:53:26 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8;
  wire n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
    n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
    n38;
  assign n10 = ~i0 & i1;
  assign n11 = ~i2 & n10;
  assign n12 = ~i3 & n11;
  assign n13 = i5 & n12;
  assign n14 = i6 & n13;
  assign n15 = ~i0 & ~i1;
  assign n16 = ~i2 & n15;
  assign n17 = ~i3 & n16;
  assign n18 = i4 & n17;
  assign n19 = i5 & n18;
  assign n20 = i0 & ~i1;
  assign n21 = ~i2 & n20;
  assign n22 = ~i3 & n21;
  assign n23 = i5 & n22;
  assign n24 = i6 & n23;
  assign n25 = ~i1 & ~i2;
  assign n26 = ~i3 & n25;
  assign n27 = i4 & n26;
  assign n28 = i6 & n27;
  assign n29 = i6 & n26;
  assign n30 = i6 & i7;
  assign n31 = i5 & n30;
  assign n32 = i4 & n31;
  assign n33 = i7 & ~n32;
  assign n34 = ~n14 & n33;
  assign n35 = ~n19 & n34;
  assign n36 = ~n24 & n35;
  assign n37 = ~n28 & n36;
  assign n38 = ~n29 & n37;
  assign i8 = n17 | ~n38;
endmodule


