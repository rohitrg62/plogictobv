// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:27:09 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8, i9, i10, i11  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8, i9, i10, i11;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
    n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
    n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n55,
    n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n182, n183,
    n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
    n316, n317;
  assign n13 = ~i0 & i1;
  assign n14 = ~i2 & n13;
  assign n15 = ~i3 & n14;
  assign n16 = ~i4 & n15;
  assign n17 = i5 & n16;
  assign n18 = i7 & n17;
  assign n19 = i0 & ~i2;
  assign n20 = ~i3 & n19;
  assign n21 = ~i4 & n20;
  assign n22 = ~i5 & n21;
  assign n23 = ~i7 & n22;
  assign n24 = i4 & n15;
  assign n25 = ~i5 & n24;
  assign n26 = i7 & n25;
  assign n27 = i0 & ~i1;
  assign n28 = ~i2 & n27;
  assign n29 = ~i3 & n28;
  assign n30 = i4 & n29;
  assign n31 = i7 & n30;
  assign n32 = i5 & n24;
  assign n33 = i7 & n32;
  assign n34 = i4 & n20;
  assign n35 = i5 & n34;
  assign n36 = i7 & n35;
  assign n37 = i1 & ~i2;
  assign n38 = ~i3 & n37;
  assign n39 = ~i4 & n38;
  assign n40 = ~i5 & n39;
  assign n41 = ~i7 & n40;
  assign n42 = ~i0 & ~i1;
  assign n43 = ~i2 & n42;
  assign n44 = i3 & n43;
  assign n45 = ~i4 & n44;
  assign n46 = ~i5 & n45;
  assign n47 = ~i7 & n46;
  assign n48 = ~n18 & ~n23;
  assign n49 = ~n26 & n48;
  assign n50 = ~n31 & n49;
  assign n51 = ~n33 & n50;
  assign n52 = ~n36 & n51;
  assign n53 = ~n41 & n52;
  assign i8 = ~n47 & n53;
  assign n55 = i4 & n44;
  assign n56 = i5 & n55;
  assign n57 = i7 & n56;
  assign n58 = i8 & n57;
  assign n59 = ~i4 & n29;
  assign n60 = i5 & n59;
  assign n61 = i7 & n60;
  assign n62 = i8 & n61;
  assign n63 = ~i1 & ~i6;
  assign n64 = ~i1 & i6;
  assign n65 = ~n63 & ~n64;
  assign n66 = i1 & ~i5;
  assign n67 = i0 & n66;
  assign n68 = ~i7 & n67;
  assign n69 = n65 & ~n68;
  assign n70 = i1 & i5;
  assign n71 = n69 & ~n70;
  assign n72 = ~n58 & ~n71;
  assign i9 = ~n62 & n72;
  assign n74 = i6 & n60;
  assign n75 = i8 & n74;
  assign n76 = i9 & n75;
  assign n77 = i2 & n42;
  assign n78 = ~i3 & n77;
  assign n79 = ~i6 & n78;
  assign n80 = i7 & n79;
  assign n81 = i8 & n80;
  assign n82 = i4 & n78;
  assign n83 = i5 & n82;
  assign n84 = i6 & n83;
  assign n85 = i8 & n84;
  assign n86 = i9 & n85;
  assign n87 = ~i4 & n14;
  assign n88 = i5 & n87;
  assign n89 = i6 & n88;
  assign n90 = ~i7 & n89;
  assign n91 = i8 & n90;
  assign n92 = i9 & n91;
  assign n93 = ~i4 & n37;
  assign n94 = ~i5 & n93;
  assign n95 = ~i6 & n94;
  assign n96 = ~i7 & n95;
  assign n97 = ~i4 & n19;
  assign n98 = ~i5 & n97;
  assign n99 = ~i6 & n98;
  assign n100 = ~i7 & n99;
  assign n101 = ~i3 & n13;
  assign n102 = i4 & n101;
  assign n103 = ~i5 & n102;
  assign n104 = i6 & n103;
  assign n105 = i7 & n104;
  assign n106 = i8 & n105;
  assign n107 = i6 & n20;
  assign n108 = ~i7 & n107;
  assign n109 = i8 & n108;
  assign n110 = ~i3 & n27;
  assign n111 = i4 & n110;
  assign n112 = ~i5 & n111;
  assign n113 = ~i6 & n112;
  assign n114 = i7 & n113;
  assign n115 = i8 & n114;
  assign n116 = i6 & n78;
  assign n117 = i7 & n116;
  assign n118 = i8 & n117;
  assign n119 = i6 & n44;
  assign n120 = ~i7 & n119;
  assign n121 = i8 & n120;
  assign n122 = i6 & n112;
  assign n123 = i7 & n122;
  assign n124 = i8 & n123;
  assign n125 = ~i4 & n28;
  assign n126 = i5 & n125;
  assign n127 = i6 & n126;
  assign n128 = ~i7 & n127;
  assign n129 = i8 & n128;
  assign n130 = i9 & n129;
  assign n131 = ~i6 & n103;
  assign n132 = i7 & n131;
  assign n133 = i8 & n132;
  assign n134 = ~i6 & ~i8;
  assign n135 = ~i7 & n134;
  assign n136 = i2 & n135;
  assign n137 = i3 & n136;
  assign n138 = i7 & n134;
  assign n139 = ~i9 & n138;
  assign n140 = ~i5 & n139;
  assign n141 = i4 & n140;
  assign n142 = ~n137 & ~n141;
  assign n143 = i9 & n138;
  assign n144 = n142 & ~n143;
  assign n145 = ~i6 & i8;
  assign n146 = ~i2 & n145;
  assign n147 = n144 & ~n146;
  assign n148 = i2 & n145;
  assign n149 = i5 & n148;
  assign n150 = i9 & n149;
  assign n151 = n147 & ~n150;
  assign n152 = i6 & ~i7;
  assign n153 = ~i4 & n152;
  assign n154 = n151 & ~n153;
  assign n155 = i4 & n152;
  assign n156 = ~i8 & n155;
  assign n157 = n154 & ~n156;
  assign n158 = i8 & n155;
  assign n159 = i2 & n158;
  assign n160 = n157 & ~n159;
  assign n161 = i6 & i7;
  assign n162 = i2 & n161;
  assign n163 = ~i5 & n162;
  assign n164 = n160 & ~n163;
  assign n165 = i5 & n162;
  assign n166 = ~i8 & n165;
  assign n167 = n164 & ~n166;
  assign n168 = ~n76 & ~n167;
  assign n169 = ~n81 & ~n168;
  assign n170 = ~n86 & ~n169;
  assign n171 = ~n92 & n170;
  assign n172 = ~n96 & n171;
  assign n173 = ~n100 & n172;
  assign n174 = ~n106 & n173;
  assign n175 = ~n109 & n174;
  assign n176 = ~n115 & ~n175;
  assign n177 = ~n118 & ~n176;
  assign n178 = ~n121 & n177;
  assign n179 = ~n124 & n178;
  assign n180 = ~n130 & n179;
  assign i11 = n133 | n180;
  assign n182 = ~i6 & n82;
  assign n183 = i8 & n182;
  assign n184 = ~i11 & n183;
  assign n185 = n32 & i9;
  assign n186 = i5 & n30;
  assign n187 = i9 & n186;
  assign n188 = ~i5 & n59;
  assign n189 = i5 & n44;
  assign n190 = i7 & n189;
  assign n191 = i8 & n190;
  assign n192 = i9 & n191;
  assign n193 = i7 & n55;
  assign n194 = i8 & n193;
  assign n195 = i4 & n14;
  assign n196 = i5 & n195;
  assign n197 = i7 & n196;
  assign n198 = i8 & n197;
  assign n199 = i9 & n198;
  assign n200 = i4 & n28;
  assign n201 = i5 & n200;
  assign n202 = i7 & n201;
  assign n203 = i8 & n202;
  assign n204 = i9 & n203;
  assign n205 = ~i5 & n16;
  assign n206 = i7 & n34;
  assign n207 = i8 & n206;
  assign n208 = n59 & ~i9;
  assign n209 = i5 & n20;
  assign n210 = i7 & n209;
  assign n211 = i8 & n210;
  assign n212 = i9 & n211;
  assign n213 = ~i7 & n98;
  assign n214 = i8 & n213;
  assign n215 = i9 & n214;
  assign n216 = n22 & i9;
  assign n217 = ~i5 & n87;
  assign n218 = ~i7 & n217;
  assign n219 = i8 & n218;
  assign n220 = ~i4 & n101;
  assign n221 = ~i5 & n220;
  assign n222 = ~i6 & n221;
  assign n223 = i7 & n222;
  assign n224 = i8 & n223;
  assign n225 = ~i11 & n224;
  assign n226 = i5 & n102;
  assign n227 = i6 & n226;
  assign n228 = i8 & n227;
  assign n229 = i9 & n228;
  assign n230 = i11 & n229;
  assign n231 = ~i4 & n110;
  assign n232 = ~i5 & n231;
  assign n233 = i6 & n232;
  assign n234 = i7 & n233;
  assign n235 = i8 & n234;
  assign n236 = i11 & n235;
  assign n237 = i6 & n221;
  assign n238 = i7 & n237;
  assign n239 = i8 & n238;
  assign n240 = i11 & n239;
  assign n241 = ~i6 & n232;
  assign n242 = i7 & n241;
  assign n243 = i8 & n242;
  assign n244 = ~i11 & n243;
  assign n245 = i4 & n77;
  assign n246 = i6 & n245;
  assign n247 = i7 & n246;
  assign n248 = i8 & n247;
  assign n249 = i11 & n248;
  assign n250 = i6 & n82;
  assign n251 = i8 & n250;
  assign n252 = i11 & n251;
  assign n253 = i5 & n19;
  assign n254 = i6 & n253;
  assign n255 = i8 & n254;
  assign n256 = i9 & n255;
  assign n257 = i11 & n256;
  assign n258 = ~i6 & n245;
  assign n259 = i7 & n258;
  assign n260 = i8 & n259;
  assign n261 = ~i11 & n260;
  assign n262 = i0 & ~i3;
  assign n263 = i4 & n262;
  assign n264 = i6 & n263;
  assign n265 = i7 & n264;
  assign n266 = i8 & n265;
  assign n267 = i11 & n266;
  assign n268 = i5 & n111;
  assign n269 = i6 & n268;
  assign n270 = i8 & n269;
  assign n271 = i9 & n270;
  assign n272 = i11 & n271;
  assign n273 = i5 & n78;
  assign n274 = i6 & n273;
  assign n275 = i8 & n274;
  assign n276 = i9 & n275;
  assign n277 = i11 & n276;
  assign n278 = ~i0 & ~i2;
  assign n279 = ~i0 & i2;
  assign n280 = ~n278 & ~n279;
  assign n281 = i0 & ~i4;
  assign n282 = n280 & ~n281;
  assign n283 = i0 & i4;
  assign n284 = ~i6 & n283;
  assign n285 = ~i11 & n284;
  assign n286 = i5 & n285;
  assign n287 = n282 & ~n286;
  assign n288 = i11 & n284;
  assign n289 = n287 & ~n288;
  assign n290 = i6 & n283;
  assign n291 = n289 & ~n290;
  assign n292 = ~n184 & ~n291;
  assign n293 = ~n185 & n292;
  assign n294 = ~n187 & n293;
  assign n295 = ~n188 & n294;
  assign n296 = ~n192 & n295;
  assign n297 = ~n194 & n296;
  assign n298 = ~n199 & n297;
  assign n299 = ~n204 & n298;
  assign n300 = ~n205 & n299;
  assign n301 = ~n207 & n300;
  assign n302 = ~n208 & n301;
  assign n303 = ~n212 & n302;
  assign n304 = ~n215 & n303;
  assign n305 = ~n216 & n304;
  assign n306 = ~n219 & n305;
  assign n307 = ~n225 & n306;
  assign n308 = ~n230 & n307;
  assign n309 = ~n236 & n308;
  assign n310 = ~n240 & n309;
  assign n311 = ~n244 & n310;
  assign n312 = ~n249 & n311;
  assign n313 = ~n252 & n312;
  assign n314 = ~n257 & n313;
  assign n315 = ~n261 & n314;
  assign n316 = ~n267 & n315;
  assign n317 = ~n272 & n316;
  assign i10 = ~n277 & n317;
endmodule


