// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:27:58 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8, i9, i10, i11  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8, i9, i10, i11;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
    n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n38, n39, n40, n41,
    n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
    n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275;
  assign n13 = i0 & ~i1;
  assign n14 = i2 & n13;
  assign n15 = ~i3 & n14;
  assign n16 = i4 & n15;
  assign n17 = i5 & n16;
  assign n18 = ~i6 & n17;
  assign n19 = ~i7 & n18;
  assign n20 = i0 & i1;
  assign n21 = i2 & n20;
  assign n22 = ~i3 & n21;
  assign n23 = ~i4 & n22;
  assign n24 = ~i5 & n23;
  assign n25 = ~i6 & n24;
  assign n26 = i7 & n25;
  assign n27 = i4 & n22;
  assign n28 = i5 & n27;
  assign n29 = ~i6 & n28;
  assign n30 = ~i7 & n29;
  assign n31 = ~i6 & n16;
  assign n32 = ~i7 & n31;
  assign n33 = ~i0 & i2;
  assign n34 = ~n19 & ~n33;
  assign n35 = ~n26 & n34;
  assign n36 = ~n30 & n35;
  assign i11 = n32 | ~n36;
  assign n38 = i3 & n21;
  assign n39 = i4 & n38;
  assign n40 = ~i5 & n39;
  assign n41 = ~i6 & n40;
  assign n42 = i7 & n41;
  assign n43 = ~i11 & n42;
  assign n44 = n19 & i11;
  assign n45 = ~i6 & n27;
  assign n46 = ~i7 & n45;
  assign n47 = ~i11 & n46;
  assign n48 = n26 & i11;
  assign n49 = i5 & n15;
  assign n50 = ~i6 & n49;
  assign n51 = ~i7 & n50;
  assign n52 = ~i11 & n51;
  assign n53 = i3 & n14;
  assign n54 = ~i4 & n53;
  assign n55 = i5 & n54;
  assign n56 = ~i6 & n55;
  assign n57 = i7 & n56;
  assign n58 = ~i11 & n57;
  assign n59 = ~i0 & ~i11;
  assign n60 = i0 & ~i11;
  assign n61 = ~i1 & n60;
  assign n62 = ~n59 & ~n61;
  assign n63 = i1 & n60;
  assign n64 = n62 & ~n63;
  assign n65 = ~i4 & i11;
  assign n66 = n64 & ~n65;
  assign n67 = i4 & i11;
  assign n68 = ~i5 & n67;
  assign n69 = n66 & ~n68;
  assign n70 = i5 & n67;
  assign n71 = n69 & ~n70;
  assign n72 = ~n43 & ~n71;
  assign n73 = ~n44 & n72;
  assign n74 = ~n47 & n73;
  assign n75 = ~n48 & n74;
  assign n76 = ~n52 & n75;
  assign i10 = ~n58 & n76;
  assign n78 = n42 & ~i10;
  assign n79 = ~i11 & n78;
  assign n80 = n46 & ~i10;
  assign n81 = ~i11 & n80;
  assign n82 = ~i0 & i1;
  assign n83 = i2 & n82;
  assign n84 = i3 & n83;
  assign n85 = ~i4 & n84;
  assign n86 = i5 & n85;
  assign n87 = ~i6 & n86;
  assign n88 = i7 & n87;
  assign n89 = i10 & n88;
  assign n90 = i11 & n89;
  assign n91 = i1 & i2;
  assign n92 = i3 & n91;
  assign n93 = ~i4 & n92;
  assign n94 = ~i6 & n93;
  assign n95 = i7 & n94;
  assign n96 = i10 & n95;
  assign n97 = i11 & n96;
  assign n98 = n30 & i11;
  assign n99 = i0 & i2;
  assign n100 = ~i3 & n99;
  assign n101 = i5 & n100;
  assign n102 = ~i6 & n101;
  assign n103 = ~i7 & n102;
  assign n104 = ~i10 & n103;
  assign n105 = ~i11 & n104;
  assign n106 = ~i0 & ~i1;
  assign n107 = i2 & n106;
  assign n108 = ~i3 & n107;
  assign n109 = ~i4 & n108;
  assign n110 = i5 & n109;
  assign n111 = ~i6 & n110;
  assign n112 = ~i7 & n111;
  assign n113 = i10 & n112;
  assign n114 = i11 & n113;
  assign n115 = i4 & n53;
  assign n116 = i5 & n115;
  assign n117 = ~i6 & n116;
  assign n118 = ~i7 & n117;
  assign n119 = i10 & n118;
  assign n120 = ~i11 & n119;
  assign n121 = i3 & n107;
  assign n122 = ~i4 & n121;
  assign n123 = ~i5 & n122;
  assign n124 = ~i6 & n123;
  assign n125 = i7 & n124;
  assign n126 = i10 & n125;
  assign n127 = i11 & n126;
  assign n128 = ~i4 & n38;
  assign n129 = ~i5 & n128;
  assign n130 = ~i6 & n129;
  assign n131 = i7 & n130;
  assign n132 = i10 & n131;
  assign n133 = ~i11 & n132;
  assign n134 = i4 & n108;
  assign n135 = ~i5 & n134;
  assign n136 = ~i6 & n135;
  assign n137 = ~i7 & n136;
  assign n138 = i10 & n137;
  assign n139 = i11 & n138;
  assign n140 = i3 & n99;
  assign n141 = ~i4 & n140;
  assign n142 = i5 & n141;
  assign n143 = ~i6 & n142;
  assign n144 = i7 & n143;
  assign n145 = ~i10 & n144;
  assign n146 = ~i11 & n145;
  assign n147 = i5 & n128;
  assign n148 = ~i6 & n147;
  assign n149 = i7 & n148;
  assign n150 = i10 & n149;
  assign n151 = ~i11 & n150;
  assign n152 = ~i6 & n54;
  assign n153 = i7 & n152;
  assign n154 = i10 & n153;
  assign n155 = ~i11 & n154;
  assign n156 = ~i3 & n83;
  assign n157 = i4 & n156;
  assign n158 = ~i6 & n157;
  assign n159 = ~i7 & n158;
  assign n160 = i10 & n159;
  assign n161 = i11 & n160;
  assign n162 = ~i0 & ~i10;
  assign n163 = i2 & n162;
  assign n164 = i1 & n163;
  assign n165 = ~i0 & i10;
  assign n166 = ~i7 & n165;
  assign n167 = ~n164 & ~n166;
  assign n168 = i0 & ~i6;
  assign n169 = n167 & ~n168;
  assign n170 = i0 & i6;
  assign n171 = ~i4 & n170;
  assign n172 = n169 & ~n171;
  assign n173 = i4 & n170;
  assign n174 = n172 & ~n173;
  assign n175 = ~n79 & ~n174;
  assign n176 = ~n81 & n175;
  assign n177 = ~n90 & ~n176;
  assign n178 = ~n97 & n177;
  assign n179 = ~n98 & n178;
  assign n180 = ~n105 & ~n179;
  assign n181 = ~n114 & n180;
  assign n182 = ~n120 & n181;
  assign n183 = ~n127 & ~n182;
  assign n184 = ~n133 & ~n183;
  assign n185 = ~n139 & n184;
  assign n186 = ~n146 & n185;
  assign n187 = ~n151 & n186;
  assign n188 = ~n155 & n187;
  assign i9 = ~n161 & n188;
  assign n190 = ~i2 & n82;
  assign n191 = i3 & n190;
  assign n192 = ~i4 & n191;
  assign n193 = ~i5 & n192;
  assign n194 = ~i6 & n193;
  assign n195 = i7 & n194;
  assign n196 = ~i9 & n195;
  assign n197 = i10 & n196;
  assign n198 = ~i11 & n197;
  assign n199 = ~i6 & n100;
  assign n200 = ~i7 & n199;
  assign n201 = i9 & n200;
  assign n202 = ~i10 & n201;
  assign n203 = i11 & n202;
  assign n204 = ~i6 & n85;
  assign n205 = i9 & n204;
  assign n206 = i10 & n205;
  assign n207 = i11 & n206;
  assign n208 = ~i6 & n99;
  assign n209 = ~i7 & n208;
  assign n210 = ~i9 & n209;
  assign n211 = ~i10 & n210;
  assign n212 = ~i11 & n211;
  assign n213 = ~i5 & n38;
  assign n214 = ~i6 & n213;
  assign n215 = ~i9 & n214;
  assign n216 = ~i10 & n215;
  assign n217 = ~i11 & n216;
  assign n218 = ~i6 & n15;
  assign n219 = ~i7 & n218;
  assign n220 = i9 & n219;
  assign n221 = i10 & n220;
  assign n222 = i11 & n221;
  assign n223 = n124 & i9;
  assign n224 = i10 & n223;
  assign n225 = i11 & n224;
  assign n226 = ~i6 & n141;
  assign n227 = ~i9 & n226;
  assign n228 = ~i10 & n227;
  assign n229 = ~i11 & n228;
  assign n230 = ~i2 & ~i6;
  assign n231 = ~i11 & n230;
  assign n232 = ~i9 & n231;
  assign n233 = i4 & n232;
  assign n234 = ~i1 & n233;
  assign n235 = i1 & n233;
  assign n236 = i7 & n235;
  assign n237 = ~n234 & ~n236;
  assign n238 = i9 & n231;
  assign n239 = n237 & ~n238;
  assign n240 = i11 & n230;
  assign n241 = n239 & ~n240;
  assign n242 = i2 & ~i6;
  assign n243 = ~i11 & n242;
  assign n244 = ~i3 & n243;
  assign n245 = i4 & n244;
  assign n246 = ~i7 & n245;
  assign n247 = n241 & ~n246;
  assign n248 = i3 & n243;
  assign n249 = i10 & n248;
  assign n250 = n247 & ~n249;
  assign n251 = i11 & n242;
  assign n252 = i7 & n251;
  assign n253 = ~i0 & n252;
  assign n254 = ~i3 & n253;
  assign n255 = n250 & ~n254;
  assign n256 = i3 & n253;
  assign n257 = ~i9 & n256;
  assign n258 = n255 & ~n257;
  assign n259 = i6 & i11;
  assign n260 = ~i7 & n259;
  assign n261 = ~i2 & n260;
  assign n262 = ~i3 & n261;
  assign n263 = n258 & ~n262;
  assign n264 = i3 & n261;
  assign n265 = i5 & n264;
  assign n266 = n263 & ~n265;
  assign n267 = ~n198 & n266;
  assign n268 = ~n203 & ~n267;
  assign n269 = ~n207 & n268;
  assign n270 = ~n207 & n269;
  assign n271 = ~n203 & n270;
  assign n272 = ~n212 & ~n271;
  assign n273 = ~n217 & n272;
  assign n274 = ~n222 & ~n273;
  assign n275 = ~n225 & n274;
  assign i8 = n229 | n275;
endmodule


