// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:28:19 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8, i9, i10, i11  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8, i9, i10, i11;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
    n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
    n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
    n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314;
  assign n13 = ~i0 & i1;
  assign n14 = ~i2 & n13;
  assign n15 = ~i3 & n14;
  assign n16 = i4 & n15;
  assign n17 = ~i5 & n16;
  assign n18 = ~i6 & n17;
  assign n19 = i7 & n18;
  assign n20 = i5 & n16;
  assign n21 = ~i6 & n20;
  assign n22 = i7 & n21;
  assign n23 = i0 & i1;
  assign n24 = ~i2 & n23;
  assign n25 = ~i3 & n24;
  assign n26 = i4 & n25;
  assign n27 = i6 & n26;
  assign n28 = ~i7 & n27;
  assign n29 = ~i4 & n25;
  assign n30 = i5 & n29;
  assign n31 = i6 & n30;
  assign n32 = ~i7 & n31;
  assign n33 = ~i3 & i6;
  assign n34 = ~i2 & n33;
  assign n35 = ~i7 & n34;
  assign n36 = i7 & n34;
  assign n37 = ~n35 & ~n36;
  assign n38 = ~n19 & n37;
  assign n39 = ~n22 & n38;
  assign n40 = ~n28 & ~n39;
  assign i11 = ~n32 & n40;
  assign n42 = ~i0 & ~i1;
  assign n43 = ~i2 & n42;
  assign n44 = ~i3 & n43;
  assign n45 = ~i6 & n44;
  assign n46 = i7 & n45;
  assign n47 = ~i11 & n46;
  assign n48 = i4 & n44;
  assign n49 = i5 & n48;
  assign n50 = ~i6 & n49;
  assign n51 = ~i11 & n50;
  assign n52 = n22 & i11;
  assign n53 = n19 & i11;
  assign n54 = ~i6 & i11;
  assign n55 = ~i7 & n54;
  assign n56 = i7 & n54;
  assign n57 = ~n55 & ~n56;
  assign n58 = i6 & i11;
  assign n59 = ~i0 & n58;
  assign n60 = ~i1 & n59;
  assign n61 = ~i3 & n60;
  assign n62 = n57 & ~n61;
  assign n63 = i3 & n60;
  assign n64 = i7 & n63;
  assign n65 = n62 & ~n64;
  assign n66 = i1 & n59;
  assign n67 = i7 & n66;
  assign n68 = n65 & ~n67;
  assign n69 = ~n47 & n68;
  assign n70 = ~n51 & n69;
  assign n71 = ~n52 & ~n70;
  assign i10 = ~n53 & n71;
  assign n73 = i5 & n44;
  assign n74 = ~i6 & n73;
  assign n75 = ~i10 & n74;
  assign n76 = ~i11 & n75;
  assign n77 = ~i6 & n48;
  assign n78 = ~i10 & n77;
  assign n79 = ~i11 & n78;
  assign n80 = ~i7 & n18;
  assign n81 = ~i10 & n80;
  assign n82 = ~i11 & n81;
  assign n83 = ~i7 & n21;
  assign n84 = ~i10 & n83;
  assign n85 = ~i11 & n84;
  assign n86 = i3 & n43;
  assign n87 = ~i4 & n86;
  assign n88 = i5 & n87;
  assign n89 = i6 & n88;
  assign n90 = i7 & n89;
  assign n91 = ~i10 & n90;
  assign n92 = ~i11 & n91;
  assign n93 = i3 & n14;
  assign n94 = i4 & n93;
  assign n95 = i5 & n94;
  assign n96 = i6 & n95;
  assign n97 = i7 & n96;
  assign n98 = ~i10 & n97;
  assign n99 = ~i11 & n98;
  assign n100 = i0 & ~i1;
  assign n101 = ~i2 & n100;
  assign n102 = ~i3 & n101;
  assign n103 = i4 & n102;
  assign n104 = i5 & n103;
  assign n105 = ~i6 & n104;
  assign n106 = i7 & n105;
  assign n107 = ~i10 & n106;
  assign n108 = ~i11 & n107;
  assign n109 = i4 & n86;
  assign n110 = ~i5 & n109;
  assign n111 = i6 & n110;
  assign n112 = i7 & n111;
  assign n113 = ~i10 & n112;
  assign n114 = ~i11 & n113;
  assign n115 = ~i5 & n103;
  assign n116 = ~i6 & n115;
  assign n117 = i7 & n116;
  assign n118 = ~i10 & n117;
  assign n119 = ~i11 & n118;
  assign n120 = ~i4 & n102;
  assign n121 = ~i6 & n120;
  assign n122 = i7 & n121;
  assign n123 = ~i10 & n122;
  assign n124 = ~i11 & n123;
  assign n125 = i6 & n103;
  assign n126 = ~i7 & n125;
  assign n127 = ~i10 & n126;
  assign n128 = i11 & n127;
  assign n129 = i3 & n24;
  assign n130 = i4 & n129;
  assign n131 = i5 & n130;
  assign n132 = i6 & n131;
  assign n133 = i7 & n132;
  assign n134 = ~i10 & n133;
  assign n135 = ~i11 & n134;
  assign n136 = ~i4 & n15;
  assign n137 = i5 & n136;
  assign n138 = ~i6 & n137;
  assign n139 = i7 & n138;
  assign n140 = ~i10 & n139;
  assign n141 = ~i11 & n140;
  assign n142 = ~i5 & n136;
  assign n143 = ~i6 & n142;
  assign n144 = i7 & n143;
  assign n145 = ~i10 & n144;
  assign n146 = ~i11 & n145;
  assign n147 = i3 & n101;
  assign n148 = ~i4 & n147;
  assign n149 = i6 & n148;
  assign n150 = i7 & n149;
  assign n151 = ~i10 & n150;
  assign n152 = ~i11 & n151;
  assign n153 = ~i5 & n130;
  assign n154 = i6 & n153;
  assign n155 = i7 & n154;
  assign n156 = ~i10 & n155;
  assign n157 = ~i11 & n156;
  assign n158 = i5 & n26;
  assign n159 = ~i6 & n158;
  assign n160 = i7 & n159;
  assign n161 = ~i10 & n160;
  assign n162 = ~i11 & n161;
  assign n163 = ~i5 & n26;
  assign n164 = ~i6 & n163;
  assign n165 = i7 & n164;
  assign n166 = ~i10 & n165;
  assign n167 = ~i11 & n166;
  assign n168 = ~i5 & n87;
  assign n169 = i6 & n168;
  assign n170 = i7 & n169;
  assign n171 = ~i10 & n170;
  assign n172 = ~i11 & n171;
  assign n173 = i6 & n120;
  assign n174 = ~i7 & n173;
  assign n175 = ~i10 & n174;
  assign n176 = i11 & n175;
  assign n177 = i6 & n163;
  assign n178 = i7 & n177;
  assign n179 = ~i10 & n178;
  assign n180 = i11 & n179;
  assign n181 = i6 & n142;
  assign n182 = i7 & n181;
  assign n183 = i10 & n182;
  assign n184 = i11 & n183;
  assign n185 = i6 & n137;
  assign n186 = i7 & n185;
  assign n187 = i10 & n186;
  assign n188 = i11 & n187;
  assign n189 = i6 & n158;
  assign n190 = i7 & n189;
  assign n191 = ~i10 & n190;
  assign n192 = i11 & n191;
  assign n193 = i7 & n31;
  assign n194 = ~i10 & n193;
  assign n195 = i11 & n194;
  assign n196 = ~i5 & n29;
  assign n197 = i6 & n196;
  assign n198 = i7 & n197;
  assign n199 = ~i10 & n198;
  assign n200 = i11 & n199;
  assign n201 = ~i7 & ~i11;
  assign n202 = ~i2 & n201;
  assign n203 = i6 & n202;
  assign n204 = ~i10 & n203;
  assign n205 = i10 & n203;
  assign n206 = i0 & n205;
  assign n207 = ~n204 & ~n206;
  assign n208 = ~i11 & n207;
  assign n209 = ~n76 & n208;
  assign n210 = ~n79 & n209;
  assign n211 = ~n82 & n210;
  assign n212 = ~n85 & n211;
  assign n213 = ~n92 & n212;
  assign n214 = ~n99 & n213;
  assign n215 = ~n108 & n214;
  assign n216 = ~n114 & n215;
  assign n217 = ~n119 & n216;
  assign n218 = ~n124 & n217;
  assign n219 = ~n128 & ~n218;
  assign n220 = ~n135 & ~n219;
  assign n221 = ~n141 & n220;
  assign n222 = ~n146 & n221;
  assign n223 = ~n152 & n222;
  assign n224 = ~n157 & n223;
  assign n225 = ~n162 & n224;
  assign n226 = ~n167 & n225;
  assign n227 = ~n172 & n226;
  assign n228 = ~n176 & ~n227;
  assign n229 = ~n180 & n228;
  assign n230 = ~n184 & n229;
  assign n231 = ~n188 & n230;
  assign n232 = ~n192 & n231;
  assign n233 = ~n195 & n232;
  assign i9 = ~n200 & n233;
  assign n235 = n80 & i9;
  assign n236 = i6 & n94;
  assign n237 = ~i7 & n236;
  assign n238 = i9 & n237;
  assign n239 = i6 & n87;
  assign n240 = ~i7 & n239;
  assign n241 = i9 & n240;
  assign n242 = n133 & i9;
  assign n243 = ~i10 & n242;
  assign n244 = ~i11 & n243;
  assign n245 = n150 & i9;
  assign n246 = ~i10 & n245;
  assign n247 = ~i11 & n246;
  assign n248 = n155 & i9;
  assign n249 = ~i10 & n248;
  assign n250 = ~i11 & n249;
  assign n251 = n160 & i9;
  assign n252 = ~i10 & n251;
  assign n253 = ~i11 & n252;
  assign n254 = n165 & i9;
  assign n255 = ~i10 & n254;
  assign n256 = ~i11 & n255;
  assign n257 = i2 & n100;
  assign n258 = i3 & n257;
  assign n259 = i4 & n258;
  assign n260 = ~i5 & n259;
  assign n261 = i6 & n260;
  assign n262 = i7 & n261;
  assign n263 = ~i9 & n262;
  assign n264 = ~i10 & n263;
  assign n265 = ~i11 & n264;
  assign n266 = n178 & ~i9;
  assign n267 = ~i10 & n266;
  assign n268 = i11 & n267;
  assign n269 = n32 & ~i10;
  assign n270 = ~i11 & n269;
  assign n271 = n19 & i9;
  assign n272 = i11 & n271;
  assign n273 = i6 & n17;
  assign n274 = i7 & n273;
  assign n275 = i9 & n274;
  assign n276 = i10 & n275;
  assign n277 = i11 & n276;
  assign n278 = ~i0 & ~i10;
  assign n279 = ~i0 & i10;
  assign n280 = ~n278 & ~n279;
  assign n281 = i0 & ~i10;
  assign n282 = ~i3 & n281;
  assign n283 = i4 & n282;
  assign n284 = ~i7 & n283;
  assign n285 = n280 & ~n284;
  assign n286 = i7 & n283;
  assign n287 = n285 & ~n286;
  assign n288 = i3 & n281;
  assign n289 = ~i2 & n288;
  assign n290 = ~i9 & n289;
  assign n291 = n287 & ~n290;
  assign n292 = i9 & n289;
  assign n293 = ~i6 & n292;
  assign n294 = ~i5 & n293;
  assign n295 = n291 & ~n294;
  assign n296 = i0 & i10;
  assign n297 = ~i7 & n296;
  assign n298 = i6 & n297;
  assign n299 = n295 & ~n298;
  assign n300 = i7 & n296;
  assign n301 = n299 & ~n300;
  assign n302 = ~n235 & ~n301;
  assign n303 = ~n238 & n302;
  assign n304 = ~n241 & n303;
  assign n305 = ~n244 & n304;
  assign n306 = ~n247 & n305;
  assign n307 = ~n250 & n306;
  assign n308 = ~n253 & n307;
  assign n309 = ~n256 & n308;
  assign n310 = ~n265 & ~n309;
  assign n311 = ~n268 & ~n310;
  assign n312 = ~n270 & ~n311;
  assign n313 = ~n184 & ~n312;
  assign n314 = ~n272 & n313;
  assign i8 = ~n277 & n314;
endmodule


