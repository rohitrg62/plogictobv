// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:26:50 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3,
    i4, i5, i6, i7  );
  input  i0, i1, i2, i3;
  output i4, i5, i6, i7;
  assign i4 = ~i0;
  assign i5 = ~i2;
  assign i6 = ~i1;
  assign i7 = ~i3;
endmodule


