// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:28:07 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8, i9, i10, i11  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8, i9, i10, i11;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
    n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
    n41, n42, n43, n44, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
    n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
    n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272;
  assign n13 = ~i0 & ~i1;
  assign n14 = i2 & n13;
  assign n15 = ~i3 & n14;
  assign n16 = ~i4 & n15;
  assign n17 = i5 & n16;
  assign n18 = i6 & n17;
  assign n19 = ~i7 & n18;
  assign n20 = i0 & ~i1;
  assign n21 = i2 & n20;
  assign n22 = i3 & n21;
  assign n23 = i4 & n22;
  assign n24 = i5 & n23;
  assign n25 = i6 & n24;
  assign n26 = i7 & n25;
  assign n27 = i3 & n14;
  assign n28 = ~i4 & n27;
  assign n29 = i5 & n28;
  assign n30 = i6 & n29;
  assign n31 = i7 & n30;
  assign n32 = i1 & ~i5;
  assign n33 = ~i1 & ~i5;
  assign n34 = ~n32 & ~n33;
  assign n35 = i5 & ~i6;
  assign n36 = n34 & ~n35;
  assign n37 = i5 & i6;
  assign n38 = ~i4 & n37;
  assign n39 = n36 & ~n38;
  assign n40 = i4 & n37;
  assign n41 = i7 & n40;
  assign n42 = n39 & ~n41;
  assign n43 = ~n19 & ~n42;
  assign n44 = ~n26 & n43;
  assign i11 = ~n31 & n44;
  assign n46 = i0 & i1;
  assign n47 = ~i2 & n46;
  assign n48 = i3 & n47;
  assign n49 = i4 & n48;
  assign n50 = i5 & n49;
  assign n51 = i6 & n50;
  assign n52 = ~i7 & n51;
  assign n53 = ~i11 & n52;
  assign n54 = ~i2 & n13;
  assign n55 = i3 & n54;
  assign n56 = ~i4 & n55;
  assign n57 = i5 & n56;
  assign n58 = ~i6 & n57;
  assign n59 = i7 & n58;
  assign n60 = i11 & n59;
  assign n61 = ~i6 & ~i7;
  assign n62 = ~i4 & n61;
  assign n63 = i4 & n61;
  assign n64 = ~i3 & n63;
  assign n65 = ~n62 & ~n64;
  assign n66 = i3 & n63;
  assign n67 = ~i11 & n66;
  assign n68 = n65 & ~n67;
  assign n69 = ~i6 & i7;
  assign n70 = n68 & ~n69;
  assign n71 = ~i3 & i6;
  assign n72 = ~i2 & n71;
  assign n73 = n70 & ~n72;
  assign n74 = i2 & n71;
  assign n75 = i4 & n74;
  assign n76 = i7 & n75;
  assign n77 = n73 & ~n76;
  assign n78 = i3 & i6;
  assign n79 = ~i0 & n78;
  assign n80 = n77 & ~n79;
  assign n81 = i0 & n78;
  assign n82 = n80 & ~n81;
  assign n83 = ~n53 & ~n82;
  assign i10 = ~n60 & n83;
  assign n85 = i0 & ~i2;
  assign n86 = i3 & n85;
  assign n87 = i4 & n86;
  assign n88 = ~i5 & n87;
  assign n89 = i6 & n88;
  assign n90 = ~i7 & n89;
  assign n91 = i10 & n90;
  assign n92 = ~i2 & i3;
  assign n93 = i4 & n92;
  assign n94 = i6 & n93;
  assign n95 = ~i10 & n94;
  assign n96 = ~i4 & n48;
  assign n97 = i5 & n96;
  assign n98 = i6 & n97;
  assign n99 = ~i7 & n98;
  assign n100 = i11 & n99;
  assign n101 = ~i0 & ~i2;
  assign n102 = i3 & n101;
  assign n103 = i4 & n102;
  assign n104 = ~i5 & n103;
  assign n105 = ~i6 & n104;
  assign n106 = i7 & n105;
  assign n107 = i10 & n106;
  assign n108 = ~i4 & n92;
  assign n109 = i6 & n108;
  assign n110 = i7 & n109;
  assign n111 = i10 & n110;
  assign n112 = i11 & n111;
  assign n113 = ~i3 & n47;
  assign n114 = ~i4 & n113;
  assign n115 = i5 & n114;
  assign n116 = ~i6 & n115;
  assign n117 = i7 & n116;
  assign n118 = i10 & n117;
  assign n119 = i11 & n118;
  assign n120 = ~i4 & i10;
  assign n121 = ~i7 & n120;
  assign n122 = i10 & ~n121;
  assign n123 = i7 & n120;
  assign n124 = ~i3 & n123;
  assign n125 = i2 & n124;
  assign n126 = n122 & ~n125;
  assign n127 = i3 & n123;
  assign n128 = n126 & ~n127;
  assign n129 = i4 & i10;
  assign n130 = ~i7 & n129;
  assign n131 = ~i5 & n130;
  assign n132 = n128 & ~n131;
  assign n133 = i7 & n129;
  assign n134 = ~i6 & n133;
  assign n135 = n132 & ~n134;
  assign n136 = i6 & n133;
  assign n137 = n135 & ~n136;
  assign n138 = ~n91 & ~n137;
  assign n139 = ~n95 & ~n138;
  assign n140 = ~n100 & ~n139;
  assign n141 = ~n107 & n140;
  assign n142 = ~n112 & n141;
  assign i9 = n119 | n142;
  assign n144 = ~i0 & i2;
  assign n145 = i4 & n144;
  assign n146 = ~i5 & n145;
  assign n147 = i6 & n146;
  assign n148 = i7 & n147;
  assign n149 = i10 & n148;
  assign n150 = i1 & ~i2;
  assign n151 = i3 & n150;
  assign n152 = i4 & n151;
  assign n153 = i5 & n152;
  assign n154 = i6 & n153;
  assign n155 = ~i9 & n154;
  assign n156 = ~i11 & n155;
  assign n157 = ~i2 & n20;
  assign n158 = ~i3 & n157;
  assign n159 = i4 & n158;
  assign n160 = i5 & n159;
  assign n161 = ~i6 & n160;
  assign n162 = ~i7 & n161;
  assign n163 = ~i9 & n162;
  assign n164 = i10 & n163;
  assign n165 = ~i3 & n144;
  assign n166 = i4 & n165;
  assign n167 = ~i5 & n166;
  assign n168 = i6 & n167;
  assign n169 = ~i7 & n168;
  assign n170 = i6 & n104;
  assign n171 = i7 & n170;
  assign n172 = i9 & n171;
  assign n173 = i10 & n172;
  assign n174 = ~i5 & n92;
  assign n175 = i6 & n174;
  assign n176 = i7 & n175;
  assign n177 = i9 & n176;
  assign n178 = i10 & n177;
  assign n179 = n106 & ~i9;
  assign n180 = i10 & n179;
  assign n181 = ~i3 & n85;
  assign n182 = i4 & n181;
  assign n183 = ~i5 & n182;
  assign n184 = ~i6 & n183;
  assign n185 = i7 & n184;
  assign n186 = i9 & n185;
  assign n187 = i10 & n186;
  assign n188 = ~i4 & n181;
  assign n189 = i5 & n188;
  assign n190 = ~i6 & n189;
  assign n191 = i7 & n190;
  assign n192 = i9 & n191;
  assign n193 = i10 & n192;
  assign n194 = i11 & n193;
  assign n195 = i6 & n92;
  assign n196 = i7 & n195;
  assign n197 = i9 & n196;
  assign n198 = i10 & n197;
  assign n199 = i11 & n198;
  assign n200 = i6 & n145;
  assign n201 = i7 & n200;
  assign n202 = i10 & n201;
  assign n203 = i11 & n202;
  assign n204 = ~i1 & ~i2;
  assign n205 = i3 & n204;
  assign n206 = i4 & n205;
  assign n207 = i5 & n206;
  assign n208 = ~i6 & n207;
  assign n209 = i7 & n208;
  assign n210 = i9 & n209;
  assign n211 = i10 & n210;
  assign n212 = ~i0 & i1;
  assign n213 = ~i2 & n212;
  assign n214 = i4 & n213;
  assign n215 = i5 & n214;
  assign n216 = i6 & n215;
  assign n217 = i7 & n216;
  assign n218 = i9 & n217;
  assign n219 = i10 & n218;
  assign n220 = i11 & n219;
  assign n221 = ~i0 & ~i6;
  assign n222 = ~i5 & n221;
  assign n223 = i5 & n221;
  assign n224 = ~i9 & n223;
  assign n225 = i7 & n224;
  assign n226 = ~n222 & ~n225;
  assign n227 = ~i0 & i6;
  assign n228 = i9 & n227;
  assign n229 = ~i1 & n228;
  assign n230 = i10 & n229;
  assign n231 = ~i7 & n230;
  assign n232 = n226 & ~n231;
  assign n233 = i7 & n230;
  assign n234 = ~i3 & n233;
  assign n235 = ~i11 & n234;
  assign n236 = n232 & ~n235;
  assign n237 = i1 & n228;
  assign n238 = n236 & ~n237;
  assign n239 = i0 & ~i7;
  assign n240 = ~i10 & n239;
  assign n241 = n238 & ~n240;
  assign n242 = i10 & n239;
  assign n243 = n241 & ~n242;
  assign n244 = i0 & i7;
  assign n245 = ~i10 & n244;
  assign n246 = ~i3 & n245;
  assign n247 = n243 & ~n246;
  assign n248 = i3 & n245;
  assign n249 = i1 & n248;
  assign n250 = n247 & ~n249;
  assign n251 = i10 & n244;
  assign n252 = ~i4 & n251;
  assign n253 = ~i2 & n252;
  assign n254 = n250 & ~n253;
  assign n255 = i2 & n252;
  assign n256 = ~i6 & n255;
  assign n257 = n254 & ~n256;
  assign n258 = i4 & n251;
  assign n259 = i3 & n258;
  assign n260 = n257 & ~n259;
  assign n261 = ~n149 & ~n260;
  assign n262 = ~n156 & ~n261;
  assign n263 = ~n164 & ~n262;
  assign n264 = ~n169 & n263;
  assign n265 = ~n173 & n264;
  assign n266 = ~n178 & n265;
  assign n267 = ~n180 & n266;
  assign n268 = ~n187 & ~n267;
  assign n269 = ~n194 & ~n268;
  assign n270 = ~n199 & n269;
  assign n271 = ~n203 & n270;
  assign n272 = ~n211 & n271;
  assign i8 = ~n220 & n272;
endmodule


