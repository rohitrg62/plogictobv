// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:28:13 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3,
    i4, i5, i6, i7  );
  input  i0, i1, i2, i3;
  output i4, i5, i6, i7;
  assign i4 = 1'b1;
  assign i5 = 1'b1;
  assign i6 = 1'b1;
  assign i7 = 1'b1;
endmodule


