// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:26:36 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8, i9, i10, i11  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8, i9, i10, i11;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n25, n26, n27,
    n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
    n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
    n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
    n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n163, n164, n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288;
  assign n13 = i0 & ~i1;
  assign n14 = i2 & n13;
  assign n15 = i3 & n14;
  assign n16 = i5 & n15;
  assign n17 = i1 & ~i5;
  assign n18 = ~i1 & ~i5;
  assign n19 = ~i2 & n18;
  assign n20 = i2 & n18;
  assign n21 = ~n19 & ~n20;
  assign n22 = ~n17 & n21;
  assign n23 = ~i5 & n22;
  assign i9 = ~n16 & ~n23;
  assign n25 = ~i0 & i2;
  assign n26 = i3 & n25;
  assign n27 = ~i4 & n26;
  assign n28 = ~i5 & n27;
  assign n29 = i7 & n28;
  assign n30 = i0 & i1;
  assign n31 = i2 & n30;
  assign n32 = ~i3 & n31;
  assign n33 = ~i4 & n32;
  assign n34 = ~i5 & n33;
  assign n35 = i7 & n34;
  assign n36 = ~i0 & i1;
  assign n37 = i2 & n36;
  assign n38 = i3 & n37;
  assign n39 = i4 & n38;
  assign n40 = ~i5 & n39;
  assign n41 = i7 & n40;
  assign n42 = i4 & n15;
  assign n43 = ~i5 & n42;
  assign n44 = i7 & n43;
  assign n45 = ~i1 & i2;
  assign n46 = i3 & n45;
  assign n47 = ~i4 & n46;
  assign n48 = ~i5 & n47;
  assign n49 = i7 & n48;
  assign n50 = i7 & n42;
  assign n51 = ~i9 & n50;
  assign n52 = i5 & n27;
  assign n53 = i7 & n52;
  assign n54 = i9 & n53;
  assign n55 = i4 & n26;
  assign n56 = i5 & n55;
  assign n57 = i7 & n56;
  assign n58 = i9 & n57;
  assign n59 = i7 & n47;
  assign n60 = ~i9 & n59;
  assign n61 = ~i7 & n56;
  assign n62 = i9 & n61;
  assign n63 = i4 & n32;
  assign n64 = i5 & n63;
  assign n65 = ~i7 & n64;
  assign n66 = i9 & n65;
  assign n67 = i4 & n14;
  assign n68 = i5 & n67;
  assign n69 = ~i7 & n68;
  assign n70 = i9 & n69;
  assign n71 = ~i3 & i6;
  assign n72 = i6 & ~n71;
  assign n73 = i3 & i6;
  assign n74 = ~i0 & n73;
  assign n75 = ~i7 & n74;
  assign n76 = n72 & ~n75;
  assign n77 = i0 & n73;
  assign n78 = ~i2 & n77;
  assign n79 = n76 & ~n78;
  assign n80 = i2 & n77;
  assign n81 = ~i7 & n80;
  assign n82 = n79 & ~n81;
  assign n83 = i7 & n80;
  assign n84 = i1 & n83;
  assign n85 = i9 & n84;
  assign n86 = n82 & ~n85;
  assign n87 = ~n29 & ~n86;
  assign n88 = ~n35 & n87;
  assign n89 = ~n41 & n88;
  assign n90 = ~n44 & n89;
  assign n91 = ~n49 & n90;
  assign n92 = ~n51 & n91;
  assign n93 = ~n54 & n92;
  assign n94 = ~n58 & ~n93;
  assign n95 = ~n60 & ~n94;
  assign n96 = ~n62 & n95;
  assign n97 = ~n66 & n96;
  assign i10 = ~n70 & n97;
  assign n99 = i7 & n55;
  assign n100 = ~i10 & n99;
  assign n101 = ~i4 & n25;
  assign n102 = i5 & n101;
  assign n103 = ~i7 & n102;
  assign n104 = i9 & n103;
  assign n105 = i10 & n104;
  assign n106 = i4 & n46;
  assign n107 = i7 & n106;
  assign n108 = ~i10 & n107;
  assign n109 = ~i5 & n67;
  assign n110 = ~i7 & n109;
  assign n111 = i10 & n110;
  assign n112 = i5 & n26;
  assign n113 = i7 & n112;
  assign n114 = i9 & n113;
  assign n115 = ~i10 & n114;
  assign n116 = i9 & n56;
  assign n117 = i5 & n14;
  assign n118 = ~i7 & n117;
  assign n119 = i9 & n118;
  assign n120 = i10 & n119;
  assign n121 = ~i7 & n106;
  assign n122 = i10 & n121;
  assign n123 = ~i7 & n55;
  assign n124 = i10 & n123;
  assign n125 = i4 & n37;
  assign n126 = ~i5 & n125;
  assign n127 = ~i7 & n126;
  assign n128 = i10 & n127;
  assign n129 = i5 & n39;
  assign n130 = i9 & n129;
  assign n131 = ~i7 & n63;
  assign n132 = i10 & n131;
  assign n133 = i5 & n32;
  assign n134 = ~i7 & n133;
  assign n135 = i9 & n134;
  assign n136 = i10 & n135;
  assign n137 = ~i1 & i3;
  assign n138 = ~i5 & n137;
  assign n139 = i3 & ~n138;
  assign n140 = i5 & n137;
  assign n141 = n139 & ~n140;
  assign n142 = i1 & i3;
  assign n143 = ~i2 & n142;
  assign n144 = i6 & n143;
  assign n145 = i9 & n144;
  assign n146 = n141 & ~n145;
  assign n147 = i2 & n142;
  assign n148 = n146 & ~n147;
  assign n149 = ~n100 & ~n148;
  assign n150 = ~n105 & n149;
  assign n151 = ~n108 & n150;
  assign n152 = ~n111 & n151;
  assign n153 = ~n108 & n152;
  assign n154 = ~n115 & n153;
  assign n155 = ~n116 & ~n154;
  assign n156 = ~n120 & ~n155;
  assign n157 = ~n122 & n156;
  assign n158 = ~n124 & n157;
  assign n159 = ~n128 & n158;
  assign n160 = ~n130 & ~n159;
  assign n161 = ~n132 & ~n160;
  assign i11 = ~n136 & n161;
  assign n163 = ~i5 & n101;
  assign n164 = ~i6 & n163;
  assign n165 = ~i10 & n164;
  assign n166 = i2 & ~i3;
  assign n167 = ~i4 & n166;
  assign n168 = ~i5 & n167;
  assign n169 = ~i6 & n168;
  assign n170 = ~i10 & n169;
  assign n171 = ~i5 & n25;
  assign n172 = ~i6 & n171;
  assign n173 = ~i10 & n172;
  assign n174 = ~i11 & n173;
  assign n175 = ~i5 & n45;
  assign n176 = ~i6 & n175;
  assign n177 = ~i10 & n176;
  assign n178 = ~i11 & n177;
  assign n179 = ~i2 & n30;
  assign n180 = i3 & n179;
  assign n181 = i4 & n180;
  assign n182 = i5 & n181;
  assign n183 = ~i6 & n182;
  assign n184 = i9 & n183;
  assign n185 = i10 & n184;
  assign n186 = ~i4 & n45;
  assign n187 = ~i5 & n186;
  assign n188 = ~i6 & n187;
  assign n189 = ~i10 & n188;
  assign n190 = ~i6 & n45;
  assign n191 = ~i9 & n190;
  assign n192 = ~i10 & n191;
  assign n193 = ~i11 & n192;
  assign n194 = ~i6 & n101;
  assign n195 = ~i10 & n194;
  assign n196 = ~i11 & n195;
  assign n197 = ~i0 & i3;
  assign n198 = i4 & n197;
  assign n199 = i6 & n198;
  assign n200 = i7 & n199;
  assign n201 = ~i10 & n200;
  assign n202 = i11 & n201;
  assign n203 = i6 & n25;
  assign n204 = i7 & n203;
  assign n205 = i10 & n204;
  assign n206 = ~i4 & n179;
  assign n207 = ~i5 & n206;
  assign n208 = ~i6 & n207;
  assign n209 = i7 & n208;
  assign n210 = i10 & n209;
  assign n211 = i4 & n25;
  assign n212 = ~i6 & n211;
  assign n213 = i10 & n212;
  assign n214 = i11 & n213;
  assign n215 = ~i6 & n186;
  assign n216 = ~i9 & n215;
  assign n217 = ~i10 & n216;
  assign n218 = ~i4 & n180;
  assign n219 = ~i5 & n218;
  assign n220 = i6 & n219;
  assign n221 = ~i7 & n220;
  assign n222 = i6 & n207;
  assign n223 = i7 & n222;
  assign n224 = i10 & n223;
  assign n225 = i6 & n211;
  assign n226 = i10 & n225;
  assign n227 = i11 & n226;
  assign n228 = i5 & n198;
  assign n229 = ~i6 & n228;
  assign n230 = ~i7 & n229;
  assign n231 = i9 & n230;
  assign n232 = i10 & n231;
  assign n233 = ~i7 & n172;
  assign n234 = ~i11 & n233;
  assign n235 = ~i6 & ~i10;
  assign n236 = ~i6 & i10;
  assign n237 = ~i7 & n236;
  assign n238 = ~i11 & n237;
  assign n239 = ~n235 & ~n238;
  assign n240 = i11 & n237;
  assign n241 = i2 & n240;
  assign n242 = n239 & ~n241;
  assign n243 = i7 & n236;
  assign n244 = ~i2 & n243;
  assign n245 = ~i3 & n244;
  assign n246 = n242 & ~n245;
  assign n247 = i6 & ~i10;
  assign n248 = ~i2 & n247;
  assign n249 = ~i3 & n248;
  assign n250 = n246 & ~n249;
  assign n251 = i3 & n248;
  assign n252 = i7 & n251;
  assign n253 = i5 & n252;
  assign n254 = n250 & ~n253;
  assign n255 = i6 & i10;
  assign n256 = ~i7 & n255;
  assign n257 = ~i2 & n256;
  assign n258 = ~i1 & n257;
  assign n259 = n254 & ~n258;
  assign n260 = i1 & n257;
  assign n261 = n259 & ~n260;
  assign n262 = i7 & n255;
  assign n263 = ~i2 & n262;
  assign n264 = ~i3 & n263;
  assign n265 = i5 & n264;
  assign n266 = n261 & ~n265;
  assign n267 = i3 & n263;
  assign n268 = n266 & ~n267;
  assign n269 = i2 & n262;
  assign n270 = n268 & ~n269;
  assign n271 = ~n165 & n270;
  assign n272 = ~n170 & n271;
  assign n273 = ~n174 & n272;
  assign n274 = ~n178 & n273;
  assign n275 = ~n185 & ~n274;
  assign n276 = ~n189 & ~n275;
  assign n277 = ~n193 & n276;
  assign n278 = ~n196 & n277;
  assign n279 = ~n202 & n278;
  assign n280 = ~n205 & n279;
  assign n281 = ~n210 & ~n280;
  assign n282 = ~n214 & n281;
  assign n283 = ~n217 & ~n282;
  assign n284 = ~n221 & ~n283;
  assign n285 = ~n224 & ~n284;
  assign n286 = ~n227 & n285;
  assign n287 = ~n232 & ~n286;
  assign n288 = ~n234 & ~n287;
  assign i8 = n234 | ~n288;
endmodule


