// Benchmark "SKOLEMFORMULA" written by ABC on Mon May  4 05:26:35 2020

module SKOLEMFORMULA ( 
    i0, i1, i2, i3, i4, i5, i6, i7,
    i8, i9, i10, i11  );
  input  i0, i1, i2, i3, i4, i5, i6, i7;
  output i8, i9, i10, i11;
  wire n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
    n27, n28, n29, n30, n31, n32, n33, n35, n36, n37, n38, n39, n40, n41,
    n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
    n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
    n84, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
    n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
    n316, n317;
  assign n13 = i1 & i2;
  assign n14 = ~i4 & n13;
  assign n15 = ~i5 & n14;
  assign n16 = i6 & n15;
  assign n17 = ~i7 & n16;
  assign n18 = i0 & i2;
  assign n19 = i3 & n18;
  assign n20 = ~i4 & n19;
  assign n21 = ~i5 & n20;
  assign n22 = i6 & n21;
  assign n23 = ~i7 & n22;
  assign n24 = ~i4 & n18;
  assign n25 = ~i5 & n24;
  assign n26 = i6 & n25;
  assign n27 = ~i7 & n26;
  assign n28 = i2 & ~i4;
  assign n29 = ~i5 & n28;
  assign n30 = i6 & n29;
  assign n31 = ~i7 & n30;
  assign n32 = ~n17 & ~n23;
  assign n33 = ~n27 & n32;
  assign i11 = ~n31 & n33;
  assign n35 = ~i0 & ~i2;
  assign n36 = ~i3 & n35;
  assign n37 = ~i4 & n36;
  assign n38 = ~i5 & n37;
  assign n39 = ~i6 & n38;
  assign n40 = i7 & n39;
  assign n41 = i3 & n13;
  assign n42 = ~i4 & n41;
  assign n43 = ~i5 & n42;
  assign n44 = ~i6 & n43;
  assign n45 = i7 & n44;
  assign n46 = ~i2 & ~i3;
  assign n47 = ~i4 & n46;
  assign n48 = ~i5 & n47;
  assign n49 = ~i6 & n48;
  assign n50 = i7 & n49;
  assign n51 = i2 & i3;
  assign n52 = ~i4 & n51;
  assign n53 = ~i5 & n52;
  assign n54 = ~i6 & n53;
  assign n55 = i7 & n54;
  assign n56 = i0 & ~i1;
  assign n57 = ~i2 & n56;
  assign n58 = i3 & n57;
  assign n59 = i4 & n58;
  assign n60 = i5 & n59;
  assign n61 = i11 & n60;
  assign n62 = ~i0 & i1;
  assign n63 = ~i2 & n62;
  assign n64 = i3 & n63;
  assign n65 = i4 & n64;
  assign n66 = i5 & n65;
  assign n67 = i11 & n66;
  assign n68 = i3 & n35;
  assign n69 = i4 & n68;
  assign n70 = ~i5 & n69;
  assign n71 = i7 & n70;
  assign n72 = i11 & n71;
  assign n73 = i0 & ~i2;
  assign n74 = ~i3 & n73;
  assign n75 = i4 & n74;
  assign n76 = ~i5 & n75;
  assign n77 = i7 & n76;
  assign n78 = i11 & n77;
  assign n79 = ~n40 & ~n45;
  assign n80 = ~n50 & n79;
  assign n81 = ~n55 & n80;
  assign n82 = ~n61 & n81;
  assign n83 = ~n67 & n82;
  assign n84 = ~n72 & n83;
  assign i8 = ~n78 & n84;
  assign n86 = ~i1 & ~i2;
  assign n87 = i3 & n86;
  assign n88 = i4 & n87;
  assign n89 = i5 & n88;
  assign n90 = ~i6 & n89;
  assign n91 = ~i7 & n90;
  assign n92 = ~i8 & n91;
  assign n93 = i5 & n69;
  assign n94 = ~i6 & n93;
  assign n95 = ~i7 & n94;
  assign n96 = ~i8 & n95;
  assign n97 = i0 & i1;
  assign n98 = ~i2 & n97;
  assign n99 = ~i3 & n98;
  assign n100 = ~i4 & n99;
  assign n101 = i5 & n100;
  assign n102 = i6 & n101;
  assign n103 = i7 & n102;
  assign n104 = i8 & n103;
  assign n105 = i11 & n104;
  assign n106 = ~i4 & n68;
  assign n107 = i5 & n106;
  assign n108 = i6 & n107;
  assign n109 = i7 & n108;
  assign n110 = i8 & n109;
  assign n111 = i11 & n110;
  assign n112 = ~i6 & n101;
  assign n113 = i7 & n112;
  assign n114 = i8 & n113;
  assign n115 = i11 & n114;
  assign n116 = i4 & n19;
  assign n117 = i5 & n116;
  assign n118 = ~i6 & n117;
  assign n119 = i7 & n118;
  assign n120 = i8 & n119;
  assign n121 = i11 & n120;
  assign n122 = ~i4 & n87;
  assign n123 = i5 & n122;
  assign n124 = i6 & n123;
  assign n125 = i7 & n124;
  assign n126 = i8 & n125;
  assign n127 = i11 & n126;
  assign n128 = ~i6 & n123;
  assign n129 = i7 & n128;
  assign n130 = i8 & n129;
  assign n131 = i11 & n130;
  assign n132 = i5 & n68;
  assign n133 = ~i6 & n132;
  assign n134 = i7 & n133;
  assign n135 = ~i8 & n134;
  assign n136 = i11 & n135;
  assign n137 = ~i6 & n107;
  assign n138 = i7 & n137;
  assign n139 = i8 & n138;
  assign n140 = i11 & n139;
  assign n141 = i6 & n93;
  assign n142 = ~i7 & n141;
  assign n143 = ~i8 & n142;
  assign n144 = i11 & n143;
  assign n145 = i5 & n87;
  assign n146 = ~i6 & n145;
  assign n147 = i7 & n146;
  assign n148 = ~i8 & n147;
  assign n149 = i11 & n148;
  assign n150 = i4 & n41;
  assign n151 = i5 & n150;
  assign n152 = ~i6 & n151;
  assign n153 = i7 & n152;
  assign n154 = i8 & n153;
  assign n155 = i11 & n154;
  assign n156 = i6 & n89;
  assign n157 = ~i7 & n156;
  assign n158 = ~i8 & n157;
  assign n159 = i11 & n158;
  assign n160 = i5 & ~i6;
  assign n161 = ~i2 & n160;
  assign n162 = ~i11 & n161;
  assign n163 = i7 & n162;
  assign n164 = i5 & ~n163;
  assign n165 = i11 & n161;
  assign n166 = ~i8 & n165;
  assign n167 = n164 & ~n166;
  assign n168 = i2 & n160;
  assign n169 = ~i0 & n168;
  assign n170 = n167 & ~n169;
  assign n171 = i0 & n168;
  assign n172 = i7 & n171;
  assign n173 = n170 & ~n172;
  assign n174 = i5 & i6;
  assign n175 = n173 & ~n174;
  assign n176 = ~n92 & n175;
  assign n177 = ~n96 & n176;
  assign n178 = ~n105 & ~n177;
  assign n179 = ~n111 & n178;
  assign n180 = ~n115 & ~n179;
  assign n181 = ~n121 & ~n180;
  assign n182 = ~n127 & n181;
  assign n183 = ~n131 & ~n182;
  assign n184 = ~n136 & ~n183;
  assign n185 = ~n140 & ~n184;
  assign n186 = ~n144 & ~n185;
  assign n187 = ~n149 & n186;
  assign n188 = ~n155 & n187;
  assign i9 = ~n159 & n188;
  assign n190 = i4 & n46;
  assign n191 = ~i5 & n190;
  assign n192 = ~i6 & n191;
  assign n193 = ~i7 & n192;
  assign n194 = i2 & n97;
  assign n195 = ~i4 & n194;
  assign n196 = i5 & n195;
  assign n197 = ~i6 & n196;
  assign n198 = i7 & n197;
  assign n199 = i8 & n198;
  assign n200 = i9 & n199;
  assign n201 = i11 & n200;
  assign n202 = i7 & n101;
  assign n203 = i11 & n202;
  assign n204 = i4 & n18;
  assign n205 = ~i5 & n204;
  assign n206 = ~i6 & n205;
  assign n207 = i7 & n206;
  assign n208 = i8 & n207;
  assign n209 = i11 & n208;
  assign n210 = ~i5 & n116;
  assign n211 = ~i6 & n210;
  assign n212 = ~i7 & n211;
  assign n213 = i7 & n107;
  assign n214 = i11 & n213;
  assign n215 = i4 & n51;
  assign n216 = ~i5 & n215;
  assign n217 = ~i6 & n216;
  assign n218 = i7 & n217;
  assign n219 = i8 & n218;
  assign n220 = i11 & n219;
  assign n221 = i4 & n63;
  assign n222 = i5 & n221;
  assign n223 = i7 & n222;
  assign n224 = i8 & n223;
  assign n225 = i11 & n224;
  assign n226 = i4 & n99;
  assign n227 = i5 & n226;
  assign n228 = i7 & n227;
  assign n229 = i8 & n228;
  assign n230 = i11 & n229;
  assign n231 = i4 & n57;
  assign n232 = i5 & n231;
  assign n233 = i7 & n232;
  assign n234 = i8 & n233;
  assign n235 = i11 & n234;
  assign n236 = i7 & n89;
  assign n237 = i8 & n236;
  assign n238 = i11 & n237;
  assign n239 = ~i8 & n192;
  assign n240 = i7 & n132;
  assign n241 = ~i8 & n240;
  assign n242 = i11 & n241;
  assign n243 = i7 & n123;
  assign n244 = i11 & n243;
  assign n245 = i5 & n52;
  assign n246 = ~i6 & n245;
  assign n247 = i7 & n246;
  assign n248 = i8 & n247;
  assign n249 = i9 & n248;
  assign n250 = i11 & n249;
  assign n251 = i7 & n145;
  assign n252 = ~i8 & n251;
  assign n253 = i11 & n252;
  assign n254 = i4 & n194;
  assign n255 = i5 & n254;
  assign n256 = ~i6 & n255;
  assign n257 = i7 & n256;
  assign n258 = i8 & n257;
  assign n259 = i9 & n258;
  assign n260 = i11 & n259;
  assign n261 = i5 & n215;
  assign n262 = ~i6 & n261;
  assign n263 = i7 & n262;
  assign n264 = i8 & n263;
  assign n265 = i9 & n264;
  assign n266 = i11 & n265;
  assign n267 = ~i7 & n152;
  assign n268 = i8 & n267;
  assign n269 = i9 & n268;
  assign n270 = i11 & n269;
  assign n271 = i4 & n13;
  assign n272 = i5 & n271;
  assign n273 = ~i6 & n272;
  assign n274 = i7 & n273;
  assign n275 = i8 & n274;
  assign n276 = i9 & n275;
  assign n277 = i11 & n276;
  assign n278 = i5 & n204;
  assign n279 = ~i6 & n278;
  assign n280 = i7 & n279;
  assign n281 = i8 & n280;
  assign n282 = i9 & n281;
  assign n283 = i11 & n282;
  assign n284 = ~i4 & ~i5;
  assign n285 = ~i4 & i5;
  assign n286 = ~n284 & ~n285;
  assign n287 = i4 & ~i6;
  assign n288 = ~i5 & n287;
  assign n289 = ~i2 & n288;
  assign n290 = i0 & n289;
  assign n291 = n286 & ~n290;
  assign n292 = i2 & n288;
  assign n293 = n291 & ~n292;
  assign n294 = i5 & n287;
  assign n295 = n293 & ~n294;
  assign n296 = i4 & i6;
  assign n297 = n295 & ~n296;
  assign n298 = ~n193 & ~n297;
  assign n299 = ~n201 & n298;
  assign n300 = ~n203 & n299;
  assign n301 = ~n209 & n300;
  assign n302 = ~n212 & n301;
  assign n303 = ~n214 & n302;
  assign n304 = ~n220 & n303;
  assign n305 = ~n225 & n304;
  assign n306 = ~n230 & n305;
  assign n307 = ~n235 & n306;
  assign n308 = ~n238 & n307;
  assign n309 = ~n239 & n308;
  assign n310 = ~n242 & n309;
  assign n311 = ~n244 & n310;
  assign n312 = ~n250 & n311;
  assign n313 = ~n253 & n312;
  assign n314 = ~n260 & n313;
  assign n315 = ~n266 & n314;
  assign n316 = ~n270 & n315;
  assign n317 = ~n277 & n316;
  assign i10 = ~n283 & n317;
endmodule


